module ALU ( nx474, nx178, nx605, nx601, src1_6, nx1901, enable_div, nx216, nx94, nx136, nx506, nx504, nx2028, src2_6, src1_3, nx1639, src2_5, src1_7, nx386, nx262, src2_2, op_code_0, bit_in, nx2019, nx1641, cycle_0, cycle_1, src1_0, nx226, nx222, nx1598, nx539, nx537, nx1782, nx308, nx1819, nx1696, nx1711, nx575, src2_1, nx459, nx593, nx455, cycle_1_div, nx1763, nx1768, nx36, nx110, nx114, src1_4, src2_4, nx1698, nx338, nx236, nx1922, tmp_rem_2, tmp_rem_3, tmp_rem_0, tmp_rem_1, tmp_rem_6, tmp_rem_4, tmp_rem_5, op_code_1, src1_1, nx50, nx1724, nx244, tmp_rem_7, op_code_2, cycle_0_div, nx415, nx1890, nx433, tmp_mul_12, enable_mul, tmp_mul_10, tmp_mul_11, nx18, src2_7, nx806, src1_2, nx567, nx64, nx60, nx1776, tmp_mul_8, tmp_mul_9, nx1778, nx102, nx730, nx10, nx128, srcCy, nx290, nx812, srcAc, src2_0, nx1945, src2_3, src1_5, op_code_3, nx12, nx22, nx252, des_acc_2, des_acc_6, desCy, des_acc_5, des_acc_1, des_acc_0, des_acc_4, des_acc_3, des_acc_7 );
input nx474, nx178, nx605, nx601, src1_6, nx1901, enable_div, nx216, nx94, nx136, nx506, nx504, nx2028, src2_6, src1_3, nx1639, src2_5, src1_7, nx386, nx262, src2_2, op_code_0, bit_in, nx2019, nx1641, cycle_0, cycle_1, src1_0, nx226, nx222, nx1598, nx539, nx537, nx1782, nx308, nx1819, nx1696, nx1711, nx575, src2_1, nx459, nx593, nx455, cycle_1_div, nx1763, nx1768, nx36, nx110, nx114, src1_4, src2_4, nx1698, nx338, nx236, nx1922, tmp_rem_2, tmp_rem_3, tmp_rem_0, tmp_rem_1, tmp_rem_6, tmp_rem_4, tmp_rem_5, op_code_1, src1_1, nx50, nx1724, nx244, tmp_rem_7, op_code_2, cycle_0_div, nx415, nx1890, nx433, tmp_mul_12, enable_mul, tmp_mul_10, tmp_mul_11, nx18, src2_7, nx806, src1_2, nx567, nx64, nx60, nx1776, tmp_mul_8, tmp_mul_9, nx1778, nx102, nx730, nx10, nx128, srcCy, nx290, nx812, srcAc, src2_0, nx1945, src2_3, src1_5, op_code_3, nx12, nx22, nx252;
output des_acc_2, des_acc_6, desCy, des_acc_5, des_acc_1, des_acc_0, des_acc_4, des_acc_3, des_acc_7;
wire nx471, sub_result_0, nx776, nx901, divsrc2_1, divsrc2_0, nx784, nx786, nx338_mul, nx1543, nx1541, nx1546, nx1547, nx176, nx174, nx1611, nx603, desCy, nx550_mul, des_acc_2, nx1882, nx1880, nx1887, nx978_div, nx1685, des1_6, nx552_div, nx929, nx1866, nx1862, nx1903, nx923, nx1906, nx1868, nx926, nx1679, nx1911, nx814, nx819, nx1914, nx182, nx444_div, nx500_div, sub_result_7, nx194_mul, nx426, nx950, nx953, nx210, nx214, divsrc1_6, divsrc1_7, divsrc1_4, divsrc1_5, divsrc1_2, divsrc1_3, divsrc1_0, divsrc1_1, nx358, nx352, nx350, nx354, des1_3, nx437, nx435, nx76, nx72, nx554_div, nx1585, nx1583, nx1581, nx1743, nx1746, nx508, nx502, nx500, nx648, nx2026, nx2021, nx2023, nx642, nx1826, nx1511, nx1513, des_acc_6, nx1519, nx410_mul, nx1828, nx910_div, nx346_div, nx1824, nx1048, nx849, nx498_div, nx910, nx913, sub_result_3, nx1950, nx916, nx919, nx851, nx853, nx855, nx1630, nx1681, nx1637, nx104, nx1706, nx829, nx826, nx821, nx823, nx543, nx989, nx546, nx983, nx554_mul, nx986, nx442, nx768, nx440, nx446, nx444, nx762, nx1559, nx1557, nx168, nx162, nx1008, nx610, nx1000, mulsrc1_1, mulsrc1_0, mulsrc1_3, sub_result_6, mulsrc1_5, mulsrc1_4, mulsrc1_7, mulsrc1_6, nx882_div, nx684, nx680, nx1854, nx1172, nx1674, nx1859, nx1676, nx1671, nx1958, nx1983, nx1981, nx1986, nx1988, nx110_div, nx861, nx865, nx536_div, nx868, nx948, nx946, nx945, nx942, nx940, nx346, nx342, nx42, nx40, nx44, nx1595, nx1591, nx1593, nx120, nx1757, nx1754, mulsrc2_0, nx1750, nx533, nx531, nx536, nx535, nx2033, nx658, nx710, nx2035, sub_result_2, nx2038, nx1847, nx1521, nx1523, nx150, nx158, nx408, nx1032, des1_4, nx2045, des_acc_5, nx2040, nx2048, nx1627, nx900, nx1963, nx1623, nx907, nx904, nx1968, nx1787, nx1780, nx1629, nx1140, nx304, nx1811, nx1714, nx836, nx1718, nx832, nx270, nx579, nx572, nx570, nx378, nx374, nx376, nx370, nx372, nx458, nx590, nx454, des1_1, nx598, nx1565, nx1561, nx1563, nx1568, nx1569, nx882, nx1625, nx1765, nx887, nx1760, nx884, nx888, nx622, des_acc_1, nx2002, nx2000, nx2006, nx2004, des_acc_0, nx756, nx750, nx694, nx980, nx1668, nx1849, nx1663, nx1661, nx480_div, nx1842, nx957, nx1991, nx1994, nx1997, nx714, nx873, nx870, nx871, nx876, nx194_div, nx879, nx978, nx1618, nx502_mul, nx1614, nx1615, sub_result_5, nx974, nx238, nx330, nx334, nx1924, nx1926, nx1920, nx442_mul, des1_5, nx1653, des_acc_4, nx56, nx1657, nx524, nx1687, nx527, nx520, nx489, des_acc_3, nx487, nx484, nx1689, nx482, nx480, nx410_div, nx937, nx975, nx1603, nx936, nx240, nx464, nx1790, nx463, nx915, nx468, nx931, nx1539, nx1537, nx1730, nx1533, nx868_div, nx410, nx414, nx258_mul, nx1025, nx1028, nx1898, nx1894, nx1896, nx572_div, nx664, nx662, nx1877, nx1651, nx1873, nx1870, nx1978, nx1793, nx1976, sub_result_1, nx1974, nx1795, nx1970, nx1152, nx1803, nx1800, nx1808, nx298, nx835, nx192, nx194, nx801, nx804, nx200, nx202, nx204, nx561, des_acc_7, nx564, nx565, nx86, nx364, nx78, nx80, nx428, nx583, nx580, nx581, nx588, nx589, nx134, nx188, nx1579, nx440_mul, nx1770, nx1773, nx897, nx890, nx893, nx519, nx518, nx515, nx514, nx517, nx516, nx510, nx513, nx2043, sub_result_4, nx739, nx146, nx2013, nx2016, nx1509, nx743, nx744, nx746, nx1739, nx1839, nx998, nx1118, nx1831, des1_2, nx1837, nx1835, nx1052, nx558, nx1947, nx966, nx960, nx1943, nx1940, nx963, nx843, nx841, nx1605, nx1607, nx2031, mulsrc1_2, nx326, nx328, nx1933, nx1931, nx1935, nx1938, nx102_div, nx498, nx550, nx552, nx554, nx556, nx491, nx1733, nx494, nx495, nx1736, nx396, nx392, nx258, nx254;
assign  nx346 = ~(nx583);
assign  nx948 = ((nx950) & (~(nx937))) | ((~(nx950)) & (nx937));
assign  nx826 = ~((nx986) & (nx1008) | ~(nx986) & (nx570));
assign  nx823 = ~((cycle_0_div) & (src2_4) | ~(cycle_0_div) & (src2_2));
assign  nx821 = ~((cycle_0_div) & (src2_5) | ~(cycle_0_div) & (src2_3));
assign  nx819 = ~((cycle_0_div) & (src2_6) | ~(cycle_0_div) & (src2_4));
assign  nx942 = ~(((src1_5) & (nx806) & (nx812)) | ((tmp_rem_5) & (nx36)));
assign  nx946 = ~(nx1983);
assign  nx945 = ~((divsrc2_0) & (nx500_div));
assign  des_acc_3 = ~((nx1866) & (nx1868) & (nx1870) & (nx1887));
assign  nx868_div = ~(((nx346_div) & (nx743)) | ((nx346_div) & (nx931)) | ((nx743) & (nx931)));
assign  nx1603 = ~(((nx1605) & (~(nx974))) | ((~(nx1605)) & (nx974)));
assign  nx480_div = ~((nx915) | (divsrc2_1));
assign  nx1605 = ~((nx1607) & ((src1_6) | (src2_6)));
assign  nx487 = ~(((nx489) & (~(nx491))) | ((~(nx489)) & (nx491)));
assign  nx762 = ~((nx756) | (nx1696) | ((nx1968) & (nx1970)));
assign  nx768 = ~((src1_5) | (nx1743));
assign  nx480 = ~(nx86);
assign  nx482 = ~(((nx342) & (~(nx923))) | ((~(nx342)) & (nx923)));
assign  nx484 = ~((src1_1) & (nx72) & ((mulsrc2_0) | (nx78)));
assign  des_acc_2 = ~((nx1824) & (nx1826) & (nx1828) & (nx1849));
assign  nx710 = ~(((nx1579) & (nx1563)) | ((nx1579) & (src2_3)) | ((nx1563) & (src2_3)));
assign  nx648 = ~((nx642) | (nx1696) | ((nx1581) & (nx1668)));
assign  nx642 = ~((nx1668) | (nx1581));
assign  nx841 = ~(((src1_0) & (nx806) & (nx812)) | ((tmp_rem_0) & (nx36)));
assign  nx1733 = ~((((nx1546) | (nx326)) & (nx10)) | (nx1568));
assign  nx1736 = ~((src1_7) & ((src1_6) | (src1_5)));
assign  nx1730 = ~((((nx1537) & (nx222)) | (nx252)) & (bit_in));
assign  nx1513 = ~((~(src2_0)) | (src1_0));
assign  nx1509 = ~((nx1513) | ((src1_0) & (nx1511)));
assign  nx1511 = ~((src2_0) & (src1_0));
assign  nx940 = ((nx942) & (~(nx931))) | ((~(nx942)) & (nx931));
assign  nx1689 = ~((src1_7) | (src2_7));
assign  nx2023 = ~(((nx946) & (src1_6)) | ((nx946) & (srcCy)) | ((src1_6) & (srcCy)));
assign  nx2026 = ~(((src1_7) & (~(srcCy))) | ((~(src1_7)) & (srcCy)));
assign  nx168 = ~((nx1760) & ((op_code_0) | (nx1757)));
assign  nx2021 = ~(((nx2023) & (~(nx2026))) | ((~(nx2023)) & (nx2026)));
assign  nx843 = ~((~(nx739)) & (divsrc2_0));
assign  nx162 = ~((nx1765) & ((nx1511) | (nx1763)));
assign  des_acc_5 = ~((nx1931) & (nx1933) & (nx1935) & (nx1958));
assign  nx1533 = ~(src1_0);
assign  nx364 = ~((nx1862) | (nx1859));
assign  mulsrc1_2 = ~(nx463);
assign  nx978_div = ~(((nx980) & (~(nx158))) | ((~(nx980)) & (nx158)));
assign  nx498_div = ~((nx929) & (nx194_div) | ~(nx929) & (nx832));
assign  des_acc_0 = ~((nx1754) & (nx1770) & (nx1773));
assign  nx182 = ~(nx1674);
assign  nx188 = ~(nx1521);
assign  nx270 = ~(((nx739) & (~(nx851))) | ((~(nx739)) & (nx851)));
assign  sub_result_1 = ((nx80) & (~(nx1519))) | ((~(nx80)) & (nx1519));
assign  divsrc1_4 = ~((nx926) & ((nx919) | (divsrc2_0)));
assign  nx410 = ~(nx1835);
assign  nx1118 = ~(((src1_7) | (nx1763)) & ((nx1627) | (nx2019)) & ((nx2021) | (nx2028)));
assign  nx739 = ~((~(tmp_rem_0)) & (cycle_0_div) & (cycle_1_div) & (src2_0));
assign  nx508 = ~(nx1559);
assign  nx463 = ~((((tmp_mul_8) & (nx386)) | (nx338_mul)) & (nx581));
assign  sub_result_2 = ((nx298) & (~(nx1539))) | ((~(nx298)) & (nx1539));
assign  nx500 = ~((src1_3) & (nx72));
assign  nx502 = ~(nx1676);
assign  nx468 = ~((nx524) & (nx226) | ~(nx524) & (nx202));
assign  sub_result_3 = ((nx458) & (~(nx1557))) | ((~(nx458)) & (nx1557));
assign  sub_result_6 = ((nx836) & (~(nx1603))) | ((~(nx836)) & (nx1603));
assign  nx983 = ~((nx572_div) & (divsrc2_0));
assign  nx986 = ~(((nx134) & (~(nx975))) | ((~(nx134)) & (nx975)));
assign  nx980 = ~(((src1_7) & (nx806) & (nx812)) | ((tmp_rem_7) & (nx36)));
assign  nx868 = ~((nx1595) & ((nx1583) | (nx1657)));
assign  nx861 = ~((divsrc2_0) & (nx270));
assign  nx502_mul = ~((src1_4) & (nx42));
assign  nx865 = ((nx1025) & (nx980)) | ((nx1025) & (nx158)) | ((nx980) & (nx158));
assign  nx214 = ~((nx812) | (nx893));
assign  nx1933 = ~(((src1_6) & (nx114)) | ((src1_4) & (nx308)));
assign  nx210 = ~(((nx527) & (nx517)) | ((nx527) & (nx519)) | ((nx517) & (nx519)));
assign  nx1837 = ~(((srcCy) & (~(src1_2))) | ((~(srcCy)) & (src1_2)));
assign  nx1835 = ~(((src1_0) & (src1_1)) | ((src1_0) & (srcCy)) | ((src1_1) & (srcCy)));
assign  nx1831 = ~(((nx352) & (nx252)) | ((src2_2) & (nx244)) | ((nx414) & (nx262)));
assign  nx1938 = ~(((nx1940) & (~(nx1943))) | ((~(nx1940)) & (nx1943)));
assign  nx915 = ~(((src1_4) & (nx806) & (nx812)) | ((tmp_rem_4) & (nx36)));
assign  nx916 = ~((nx2006) | (nx910) | ((nx2000) & (nx2002)));
assign  nx913 = ~((cycle_0_div) & (src2_3) | ~(cycle_0_div) & (src2_1));
assign  nx603 = ~((nx386) & (tmp_mul_10) & (nx346));
assign  nx910 = ~((src1_5) | (src1_6) | (nx1743));
assign  nx338_mul = ~((nx579) & (nx575) | ~(nx579) & (nx572));
assign  des_acc_7 = ~((nx2013) & (nx2016) & (nx2033) & (nx2035));
assign  nx1607 = ~((src2_6) & (src1_6));
assign  divsrc2_1 = ~((nx865) | (nx134) | (nx801));
assign  nx1790 = ~((nx326) | (srcAc));
assign  nx1795 = ~(((src1_0) & (nx308)) | ((sub_result_1) & (nx94)));
assign  nx1793 = ~(((src1_2) & (nx114)) | ((divsrc1_1) & (enable_div)));
assign  mulsrc1_1 = ((nx572) & (~(nx579))) | ((~(nx572)) & (nx579));
assign  nx572_div = ~(((nx570) & (~(nx986))) | ((~(nx570)) & (nx986)));
assign  nx326 = ~(nx1854);
assign  nx328 = ~(nx1790);
assign  divsrc1_3 = ~((nx907) & ((nx901) | (divsrc2_0)));
assign  nx1765 = ~((src2_0) & ((nx136) | (nx128)));
assign  nx258_mul = ~(((nx561) & (nx552)) | ((nx561) & (nx554_mul)) | ((nx552) & (nx554_mul)));
assign  nx1760 = ~((((src1_0) & (nx128)) | (nx162)) & (op_code_0));
assign  nx558 = ~((((src1_7) & (nx72)) | (nx258_mul)) & (nx565));
assign  divsrc1_2 = ~((nx887) & ((nx879) | (divsrc2_0)));
assign  nx543 = ~(((nx254) & (~(nx550_mul)) & (~(nx539))) | ((~(nx254)) & (nx550_mul) & (~(nx539))) | ((~(nx254)) & (~(nx550_mul)) & (nx539)) | ((nx254) & (nx550_mul) & (nx539)));
assign  nx1986 = ~(((src1_6) & (~(srcCy))) | ((~(src1_6)) & (srcCy)));
assign  nx1983 = ~(((nx814) & (src1_5)) | ((nx814) & (srcCy)) | ((src1_5) & (srcCy)));
assign  nx1981 = ~(((nx1983) & (~(nx1986))) | ((~(nx1983)) & (nx1986)));
assign  nx1547 = ~(src1_1);
assign  nx1546 = ~(((nx1736) & (~(srcCy)) & (~(nx1032))) | ((~(nx1736)) & (srcCy) & (~(nx1032))) | ((~(nx1736)) & (~(srcCy)) & (nx1032)) | ((nx1736) & (srcCy) & (nx1032)));
assign  nx1543 = ~((src2_2) & (src1_2));
assign  nx1541 = ~((nx1543) & ((src1_2) | (src2_2)));
assign  nx1988 = ~(((nx870) & (nx252)) | ((src2_6) & (nx664)));
assign  nx134 = ~((cycle_1_div) & (nx989) | ~(cycle_1_div) & (nx913));
assign  sub_result_7 = ~(((nx1615) & (~(nx1627))) | ((~(nx1615)) & (nx1627)));
assign  nx428 = ~(((nx426) & (~(nx910_div))) | ((~(nx426)) & (nx910_div)));
assign  nx786 = ~(((nx776) & (~(nx784))) | ((~(nx776)) & (nx784)));
assign  nx1618 = ~((nx1614) | (nx1639));
assign  nx784 = ~((nx1854) & (nx1537) & (nx1736));
assign  des1_2 = ~((nx1831) & (nx1839));
assign  mulsrc1_6 = ~((((nx455) | (nx433)) & (nx589)) | (nx410_mul));
assign  nx426 = ~((nx890) & (nx214) | ~(nx890) & (nx835));
assign  nx304 = ~((nx543) & (nx539) | ~(nx543) & (nx468));
assign  nx192 = ~((nx812) | (nx823));
assign  nx1870 = ~(((des1_3) & (nx564)) | ((sub_result_3) & (nx94)));
assign  nx1873 = ~(((nx502) & (nx252)) | ((src2_3) & (nx244)) | ((nx554) & (nx262)));
assign  nx1877 = ~(((nx410) & (srcCy)) | ((nx410) & (src1_2)) | ((srcCy) & (src1_2)));
assign  nx410_mul = ~(nx598);
assign  nx1826 = ~(((src1_3) & (nx114)) | ((src1_1) & (nx308)));
assign  nx258 = ~(((src1_0) & (~(nx1808))) | ((~(src1_0)) & (nx1808)));
assign  mulsrc2_0 = (src1_0) & (nx42);
assign  nx1978 = ~(((des1_6) & (nx290)) | ((sub_result_6) & (nx94)));
assign  nx550 = ~(nx1877);
assign  nx1970 = ~(((nx1583) & (~(nx1593))) | ((~(nx1583)) & (nx1593)));
assign  nx254 = ~(((nx546) & (nx533)) | ((nx546) & (nx535)) | ((nx533) & (nx535)));
assign  nx1976 = ~(((src1_7) & (nx114)) | ((src1_5) & (nx308)));
assign  divsrc1_0 = ~((((divsrc2_0) & (nx238)) | (nx841)) & (nx843));
assign  nx1974 = ~(((mulsrc1_6) & (enable_mul)) | ((divsrc1_6) & (enable_div)));
assign  nx957 = ~((nx552_div) | ((divsrc2_1) & (nx554_div)));
assign  nx814 = ~(nx1940);
assign  nx950 = ~((nx174) | ((cycle_0_div) & (src2_1) & (nx812)));
assign  nx953 = ~(((src1_6) & (nx806) & (nx812)) | ((tmp_rem_6) & (nx36)));
assign  nx1887 = ~((nx520) | ((nx1854) & (srcAc) & (nx494)));
assign  nx1882 = ~((nx536) | ((src1_3) & (nx216)) | ((nx508) & (nx222)));
assign  nx1803 = ~(((nx182) & (nx252)) | ((src2_1) & (nx244)) | ((nx258) & (nx262)));
assign  nx1800 = ~((nx200) | ((des1_1) & (nx290)));
assign  nx1808 = ~(((src1_1) & (~(srcCy))) | ((~(src1_1)) & (srcCy)));
assign  nx1569 = ((nx580) & (~(nx710))) | ((~(nx580)) & (nx710));
assign  nx1757 = ~(((nx1533) & (op_code_1) & (op_code_2)) | ((nx40) & (nx128)));
assign  nx1750 = ~((nx110) & (src1_0) & (nx1698));
assign  nx776 = ~((nx1963) & ((src1_5) | (nx768)));
assign  nx1968 = ~(nx642);
assign  nx552_div = ~((nx953) | (divsrc2_1));
assign  nx78 = ~(nx444);
assign  nx500_div = ~(((nx498_div) & (~(nx948))) | ((~(nx498_div)) & (nx948)));
assign  nx76 = ~((((nx1776) & (nx1778)) | (nx1533)) & (nx1780));
assign  nx756 = ~((nx1970) | (nx1968));
assign  nx1052 = ~((nx2040) & ((nx1768) | (nx2038)));
assign  nx72 = (src2_7) & ~(cycle_0) & ~(cycle_1) | (src2_5) & (cycle_0) & ~(cycle_1) | (src2_3) & ~(cycle_0) & (cycle_1) | (src2_1) & (cycle_0) & (cycle_1);
assign  nx580 = ~((~(nx458)) & (nx1557));
assign  nx579 = ~(((nx565) & (~(nx575))) | ((~(nx565)) & (nx575)));
assign  nx581 = ~((nx386) & (tmp_mul_8) & (nx338_mul));
assign  nx583 = ~((~(nx581)) & (nx386) & (tmp_mul_9));
assign  nx102_div = ~((((src2_5) | (src2_6)) & (nx806)) | (src2_7));
assign  nx588 = ~((nx980) | (divsrc2_1));
assign  nx298 = ~((~(nx80)) & (nx1519));
assign  nx440_mul = ~(((nx442_mul) & (~(nx444))) | ((~(nx442_mul)) & (nx444)));
assign  nx2013 = ~((nx1152) & (nx50));
assign  nx2016 = ~((op_code_0) & (nx1140) | ~(op_code_0) & (nx1118));
assign  nx174 = ~((nx812) | (nx821));
assign  nx176 = ~(nx950);
assign  nx1615 = ~(((nx978) & (~(nx1623))) | ((~(nx978)) & (nx1623)));
assign  nx1614 = ~(((nx1637) & (src2_7)) | ((nx1637) & (nx1615)) | ((src2_7) & (nx1615)));
assign  nx1611 = ~(src1_5);
assign  nx378 = ~(nx589);
assign  nx1593 = ~((nx1595) & ((src1_5) | (src2_5)));
assign  nx376 = (nx1746) | ((src1_1) & (src1_2));
assign  nx1595 = ~((src2_5) & (src1_5));
assign  nx374 = ~(nx603);
assign  nx372 = ~((nx998) | ((divsrc2_1) & (nx238)));
assign  nx1591 = ((nx1593) & (~(nx1585))) | ((~(nx1593)) & (nx1585));
assign  nx370 = ~((nx364) | (nx1696) | ((nx1859) & (nx1862)));
assign  nx194 = ~((nx1685) | (nx1687));
assign  nx1849 = ~((nx370) | ((nx376) & (nx328) & (nx338)));
assign  nx936 = ~(((nx1607) | (nx1724)) & ((src1_6) | (nx1711)));
assign  nx960 = ((nx953) & (~(nx950))) | ((~(nx953)) & (nx950));
assign  nx517 = ~((src1_4) & (nx72));
assign  nx518 = ~(((nx346_div) & (~(nx940))) | ((~(nx346_div)) & (nx940)));
assign  nx454 = ~(((nx1547) & (nx1513)) | ((nx1547) & (src2_1)) | ((nx1513) & (src2_1)));
assign  nx104 = (nx819) & (nx821) & (nx823) & (nx102_div);
assign  nx743 = ~(nx942);
assign  nx458 = ~((~(nx298)) & (nx1539));
assign  nx1539 = ~(((nx1541) & (~(nx454))) | ((~(nx1541)) & (nx454)));
assign  nx515 = ~(((nx517) & (~(nx519))) | ((~(nx517)) & (nx519)));
assign  nx516 = ~((nx942) | (divsrc2_1));
assign  nx513 = ~(nx146);
assign  nx514 = ~((nx1679) | (nx1681));
assign  nx855 = ~(nx334);
assign  nx1048 = ~((nx1778) | ((nx2043) & (nx2045)));
assign  nx851 = ((nx849) & (~(nx853))) | ((~(nx849)) & (nx853));
assign  nx849 = ~((src2_1) & (cycle_0_div) & (cycle_1_div));
assign  nx989 = ~((cycle_0_div) & (src2_7) | ~(cycle_0_div) & (src2_5));
assign  nx1947 = ~(((nx744) & (nx252)) | ((src2_5) & (nx664)));
assign  nx836 = ~((~(nx714)) & (nx1591));
assign  nx510 = ~(((nx150) & (~(nx515)) & (~(nx506))) | ((~(nx150)) & (nx515) & (~(nx506))) | ((~(nx150)) & (~(nx515)) & (nx506)) | ((nx150) & (nx515) & (nx506)));
assign  nx346_div = ~(((nx871) & (nx915)) | ((nx871) & (nx204)) | ((nx915) & (nx204)));
assign  nx1924 = ~(src1_4);
assign  nx204 = ~((nx812) | (nx913));
assign  nx1920 = ~((nx216) | ((nx1537) & (nx244)));
assign  nx202 = ~((nx510) & (nx506) | ~(nx510) & (nx471));
assign  nx200 = ~((nx194) | (nx1696) | ((nx1687) & (nx1685)));
assign  nx1842 = ~((src1_2) | (src2_2));
assign  des1_5 = ~((nx1947) & (nx1950) & ((nx1938) | (nx1945)));
assign  nx853 = ~((nx372) | ((nx855) & (divsrc2_1)));
assign  nx926 = ~((divsrc2_0) & (nx464));
assign  nx923 = ~(((nx915) & (~(nx204))) | ((~(nx915)) & (nx204)));
assign  nx194_mul = ~((nx120) & (nx480) | ~(nx120) & (nx474));
assign  nx829 = ~((nx948) & (nx950) | ~(nx948) & (nx498_div));
assign  nx998 = ~(((src1_1) & (nx806) & (nx812)) | ((tmp_rem_1) & (nx36)));
assign  nx1627 = ~((nx1629) & ((src1_7) | (src2_7)));
assign  nx1625 = ~(src2_6);
assign  nx1623 = ~(((src1_6) & (nx974)) | ((src1_6) & (nx1625)) | ((nx974) & (nx1625)));
assign  nx1152 = ((nx1651) & (~(nx1627))) | ((~(nx1651)) & (nx1627));
assign  nx1787 = ~(((mulsrc1_1) & (enable_mul)) | ((nx330) & (nx338)));
assign  nx1780 = ~((nx56) | ((nx1641) & (src1_7) & (nx1782)));
assign  nx330 = ~(((src1_1) & (~(nx1790))) | ((~(src1_1)) & (nx1790)));
assign  nx80 = ~((nx1509) & (srcCy));
assign  nx334 = ~((~(tmp_rem_1)) & (src2_0) & (cycle_0_div) & (cycle_1_div));
assign  nx1657 = ~((src1_5) | (src2_5));
assign  nx1714 = ~(nx1172);
assign  nx1651 = ((nx1653) & (~(nx882))) | ((~(nx1653)) & (nx882));
assign  nx1718 = ~((srcCy) & ((nx22) | (nx252) | (nx1598)));
assign  nx1653 = ~(((nx868) & (src1_6)) | ((nx868) & (src2_6)) | ((src1_6) & (src2_6)));
assign  nx354 = ~(((nx868_div) & (nx953)) | ((nx868_div) & (nx176)) | ((nx953) & (nx176)));
assign  nx1028 = ~(nx1739);
assign  nx1537 = ~(srcCy);
assign  sub_result_0 = ~((nx80) & ((srcCy) | (nx1509)));
assign  nx1025 = ~(nx354);
assign  nx414 = ((nx1835) & (~(nx1837))) | ((~(nx1835)) & (nx1837));
assign  nx146 = ~(((nx484) & (nx489)) | ((nx484) & (nx491)) | ((nx489) & (nx491)));
assign  nx524 = ~(((nx210) & (~(nx531)) & (~(nx537))) | ((~(nx210)) & (nx531) & (~(nx537))) | ((~(nx210)) & (~(nx531)) & (nx537)) | ((nx210) & (nx531) & (nx537)));
assign  mulsrc1_7 = ((nx598) & (~(nx605))) | ((~(nx598)) & (nx605));
assign  mulsrc1_5 = ~((((nx601) | (nx433)) & (nx603)) | (nx378));
assign  nx897 = ~(((src1_3) & (nx806) & (nx812)) | ((tmp_rem_3) & (nx36)));
assign  nx890 = ~(((nx214) & (~(nx879))) | ((~(nx214)) & (nx879)));
assign  nx893 = ~((cycle_0_div) & (src2_2) | ~(cycle_0_div) & (src2_0));
assign  des1_3 = ~((nx1873) & (nx1882));
assign  nx561 = ~(nx254);
assign  nx565 = ~((nx258_mul) & (src1_7) & (nx72));
assign  nx564 = ~((~(nx440)) & (nx1819));
assign  nx966 = ~(((nx158) & (~(nx957))) | ((~(nx158)) & (nx957)));
assign  nx963 = ~((divsrc2_0) & (nx536_div));
assign  des1_6 = ~((nx1988) & (nx1991) & ((nx1981) | (nx1945)));
assign  nx804 = ~(((nx1595) | (nx1724)) & ((src1_5) | (nx1711)));
assign  nx801 = ~((((nx110_div) | (cycle_0_div)) & (cycle_1_div)) | (nx104));
assign  nx86 = ~((nx433) | (nx415) | (nx435));
assign  nx1847 = ~((~(op_code_3)) & (op_code_0) & (nx1790) & (op_code_2));
assign  nx536_div = ((nx829) & (~(nx966))) | ((~(nx829)) & (nx966));
assign  nx1811 = ~((nx240) | ((src1_1) & (nx216)) | ((nx188) & (nx222)));
assign  nx442_mul = ~((src1_1) & (nx72));
assign  nx1743 = ~((src1_4) & (nx326));
assign  nx1746 = ~((src1_2) | (src1_1));
assign  nx1739 = ~((nx1736) & ((src1_6) | (src1_5) | (src1_7)));
assign  nx1963 = ~((~(nx1743)) & (src1_5));
assign  nx664 = (srcCy) & (nx244);
assign  nx662 = ~((nx1924) | ((nx1920) & (nx1922)));
assign  nx744 = ~(nx1657);
assign  des_acc_4 = ~((nx1894) & (nx1896) & (nx1898) & (nx1926));
assign  nx1839 = ~((nx396) | ((src1_2) & (nx216)) | ((nx358) & (nx222)));
assign  nx680 = ~(nx1906);
assign  nx589 = ~((nx386) & (tmp_mul_11) & (nx374));
assign  nx590 = ~(((nx354) & (~(nx978_div))) | ((~(nx354)) & (nx978_div)));
assign  nx598 = ~((nx386) & (tmp_mul_12) & (nx378));
assign  nx410_div = ~(((nx334) & (~(nx882_div))) | ((~(nx334)) & (nx882_div)));
assign  nx610 = ~((~(src1_4)) & (nx1854));
assign  nx556 = ~(((nx558) & (~(nx567))) | ((~(nx558)) & (nx567)));
assign  nx2006 = ~(nx784);
assign  nx2004 = ~((src1_6) | (src1_5));
assign  nx2002 = ~((nx2004) | ((src1_5) & (src1_6)));
assign  nx2000 = ~(nx768);
assign  des1_4 = ~((nx1903) & (nx1914) & ((nx1581) | (nx1901)));
assign  nx554 = ((nx1877) & (~(nx1880))) | ((~(nx1877)) & (nx1880));
assign  nx1663 = ~(nx756);
assign  nx342 = ~(((nx873) & (nx897)) | ((nx873) & (nx214)) | ((nx897) & (nx214)));
assign  nx1581 = ~((nx1585) | ((src1_4) & (nx1583)));
assign  nx1579 = ~(src1_3);
assign  des_acc_1 = ~((nx1787) & (nx1793) & (nx1795) & (nx1800));
assign  nx1926 = ~((nx648) | ((nx610) & (nx1743) & (nx338)));
assign  nx552 = ~((src1_6) & (nx72));
assign  nx56 = ~((nx44) | (nx1696) | ((nx1509) & (nx1537)));
assign  nx1940 = ~(((nx680) & (src1_4)) | ((nx680) & (srcCy)) | ((src1_4) & (srcCy)));
assign  nx464 = ((nx832) & (~(nx929))) | ((~(nx832)) & (nx929));
assign  nx1563 = ~(((src1_2) & (nx454)) | ((src1_2) & (nx1565)) | ((nx454) & (nx1565)));
assign  nx1565 = ~(src2_2);
assign  nx1559 = ~((nx1561) & ((src1_3) | (src2_3)));
assign  nx554_mul = ~((src1_7) & (nx42));
assign  nx110_div = ~((src2_7) | (src2_6));
assign  nx1568 = ~((nx1750) & ((nx60) | (bit_in) | (nx64)));
assign  nx1561 = ~((src2_3) & (src1_3));
assign  nx520 = ~((nx514) | (nx1696) | ((nx1681) & (nx1679)));
assign  nx519 = ~((src1_5) & (nx42));
assign  nx1943 = ~(((src1_5) & (~(srcCy))) | ((~(src1_5)) & (srcCy)));
assign  nx527 = ~(nx150);
assign  nx919 = ~((nx480_div) | ((divsrc2_1) & (nx482)));
assign  nx444 = ~((src1_2) & (nx42));
assign  nx446 = ((nx873) & (~(nx904))) | ((~(nx873)) & (nx904));
assign  nx440 = ~((nx1847) & ((op_code_0) | (nx12)));
assign  nx442 = ~((~(nx440)) & (nx1819));
assign  nx554_div = ((nx868_div) & (~(nx960))) | ((~(nx868_div)) & (nx960));
assign  nx882_div = ((nx884) & (~(nx849))) | ((~(nx884)) & (nx849));
assign  nx1911 = ~(((src1_4) & (~(srcCy))) | ((~(src1_4)) & (srcCy)));
assign  nx1914 = ~((((nx664) | (nx252)) & (src2_4)) | (nx662));
assign  nx238 = ~((~(src2_0)) | (nx730));
assign  nx1854 = ~((src1_3) & ((src1_2) | (src1_1)));
assign  nx835 = ~((nx851) & (nx849) | ~(nx851) & (nx739));
assign  nx937 = ~((nx516) | ((divsrc2_1) & (nx518)));
assign  nx832 = ~((nx910_div) & (nx1000) | ~(nx910_div) & (nx426));
assign  nx533 = ~((src1_5) & (nx72));
assign  nx622 = ~((nx1561) & ((nx1671) | (nx1676)));
assign  nx929 = ((nx931) & (~(nx919))) | ((~(nx931)) & (nx919));
assign  nx931 = ~((nx192) | ((cycle_0_div) & (src2_0) & (nx812)));
assign  nx550_mul = ~(((nx552) & (~(nx554_mul))) | ((~(nx552)) & (nx554_mul)));
assign  nx910_div = ~(((nx204) & (~(nx901))) | ((~(nx204)) & (nx901)));
assign  divsrc1_5 = ~((nx945) & ((nx937) | (divsrc2_0)));
assign  nx1637 = ~(src1_7);
assign  nx1880 = ~(((srcCy) & (~(src1_3))) | ((~(srcCy)) & (src1_3)));
assign  desCy = ~((nx1706) & (nx1718) & (nx1730) & (nx1733));
assign  nx1140 = ~(((nx1629) | (nx1763)) & ((nx2028) | (nx2031)) & ((nx1689) | (nx2019)));
assign  nx1630 = ~(((srcCy) | (nx1711)) & ((nx1714) | (nx1696)));
assign  nx1629 = ~((src2_7) & (src1_7));
assign  mulsrc1_0 = ~(((nx304) & (~(nx556))) | ((~(nx304)) & (nx556)));
assign  nx714 = ~((nx1581) & (nx1569));
assign  nx2040 = ~((nx1048) | ((nx1782) & (op_code_1) & (src1_6)));
assign  nx2045 = ~((nx784) & (nx2048) & ((nx910) | (nx1028)));
assign  sub_result_5 = ((nx714) & (~(nx1591))) | ((~(nx714)) & (nx1591));
assign  nx2043 = ~((nx1854) & (nx1537) & (src1_7) & (nx2004));
assign  nx495 = ~(((nx146) & (~(nx498)) & (~(nx504))) | ((~(nx146)) & (nx498) & (~(nx504))) | ((~(nx146)) & (~(nx498)) & (nx504)) | ((nx146) & (nx498) & (nx504)));
assign  nx2048 = ~(nx1032);
assign  nx491 = ~((src1_3) & (nx42));
assign  nx489 = ~((src1_2) & (nx72));
assign  nx658 = ~(nx1920);
assign  nx1706 = ~((nx1630) | (nx1618) | ((src1_7) & (nx102)));
assign  nx1032 = ~((~(nx910)) | (nx1739));
assign  nx1679 = ~(((nx1671) & (~(nx1559))) | ((~(nx1671)) & (nx1559)));
assign  nx1681 = ~(nx364);
assign  nx240 = ~(((nx1523) | (nx1724)) & ((src1_1) | (nx1711)));
assign  nx1685 = ~(((nx1511) & (~(nx1521))) | ((~(nx1511)) & (nx1521)));
assign  nx1687 = ~(nx44);
assign  nx1519 = ((nx1521) & (~(nx1513))) | ((~(nx1521)) & (nx1513));
assign  nx1521 = ~((nx1523) & ((src1_1) | (src2_1)));
assign  nx1523 = ~((src2_1) & (src1_1));
assign  nx2035 = ~((nx1052) | ((sub_result_7) & (nx94)) | ((src1_7) & (nx22)));
assign  nx2033 = ~(((mulsrc1_7) & (enable_mul)) | ((divsrc1_7) & (enable_div)));
assign  nx150 = ~(((nx513) & (nx500)) | ((nx513) & (nx502_mul)) | ((nx500) & (nx502_mul)));
assign  nx2031 = ~((srcCy) & (src2_7) | ~(srcCy) & (src1_7));
assign  nx746 = ~(nx884);
assign  nx408 = ~((nx884) | (divsrc2_1));
assign  nx158 = ~((cycle_1_div) & (nx819) | ~(cycle_1_div) & (nx893));
assign  nx2038 = ~(((src1_0) & (nx18)) | ((srcCy) & (nx1698)));
assign  mulsrc1_4 = ~((((nx459) | (nx433)) & (nx583)) | (nx374));
assign  nx396 = ~(((nx1543) | (nx1724)) & ((src1_2) | (nx1711)));
assign  nx498 = ~(((nx500) & (~(nx502_mul))) | ((~(nx500)) & (nx502_mul)));
assign  nx194_div = ~(nx931);
assign  nx1898 = ~(((des1_4) & (nx290)) | ((sub_result_4) & (nx94)));
assign  des1_1 = ~((nx1803) & (nx1811));
assign  nx1894 = ~(((mulsrc1_4) & (enable_mul)) | ((divsrc1_4) & (enable_div)));
assign  nx1896 = ~(((src1_5) & (nx114)) | ((src1_3) & (nx308)));
assign  nx1958 = ~((nx762) | ((nx338) & (nx786)));
assign  nx392 = ((nx835) & (~(nx890))) | ((~(nx835)) & (nx890));
assign  nx471 = ~((nx495) & (nx178) | ~(nx495) & (nx194_mul));
assign  divsrc1_7 = ~((nx983) & ((nx975) | (divsrc2_0)));
assign  nx570 = ~((nx966) & (nx158) | ~(nx966) & (nx829));
assign  nx572 = ~((nx556) & (nx236) | ~(nx556) & (nx304));
assign  nx975 = ~((nx588) | ((nx590) & (divsrc2_1)));
assign  nx978 = ~((~(nx836)) & (nx1603));
assign  nx1935 = ~(((des1_5) & (nx290)) | ((sub_result_5) & (nx94)));
assign  nx870 = ~(nx1994);
assign  nx871 = ~(nx342);
assign  nx873 = ~(((nx334) & (nx746)) | ((nx334) & (nx849)) | ((nx746) & (nx849)));
assign  nx876 = ~(nx1605);
assign  nx884 = ~(((src1_2) & (nx806) & (nx812)) | ((tmp_rem_2) & (nx36)));
assign  nx879 = ~((nx408) | ((divsrc2_1) & (nx410_div)));
assign  nx1824 = ~(((mulsrc1_2) & (enable_mul)) | ((divsrc1_2) & (enable_div)));
assign  nx882 = ~((nx1661) | (nx1663));
assign  nx1828 = ~(((des1_2) & (nx442)) | ((sub_result_2) & (nx94)));
assign  nx887 = ~((divsrc2_0) & (nx392));
assign  nx888 = ~((nx882) | (nx1696) | ((nx1663) & (nx1661)));
assign  nx494 = ~((nx1890) | ((nx1746) & (nx1579)));
assign  nx1770 = ~(((src1_1) & (nx114)) | ((divsrc1_0) & (enable_div)));
assign  nx1773 = ~((nx76) | ((sub_result_0) & (nx94)) | ((srcCy) & (nx102)));
assign  nx904 = ~(((nx897) & (~(nx214))) | ((~(nx897)) & (nx214)));
assign  nx900 = (nx1854) & (src1_6) & (nx1537) & (nx1736);
assign  nx901 = ~((nx444_div) | ((divsrc2_1) & (nx446)));
assign  nx750 = ~(nx1593);
assign  nx907 = ~((divsrc2_0) & (nx428));
assign  nx1661 = ((nx868) & (~(nx1605))) | ((~(nx868)) & (nx1605));
assign  nx444_div = ~((nx897) | (divsrc2_1));
assign  nx1931 = ~(((mulsrc1_5) & (enable_mul)) | ((divsrc1_5) & (enable_div)));
assign  nx1172 = ~((nx1629) & ((nx1651) | (nx1689)));
assign  nx1754 = ~((nx168) | ((mulsrc1_0) & (enable_mul)));
assign  nx1866 = ~(((mulsrc1_3) & (enable_mul)) | ((divsrc1_3) & (enable_div)));
assign  mulsrc1_3 = ~((((nx593) | (nx433)) & (nx581)) | (nx346));
assign  nx1668 = ~(((nx622) & (~(nx514))) | ((~(nx622)) & (nx514)));
assign  nx350 = ~((nx1523) & ((nx1511) | (nx1674)));
assign  nx352 = ~(nx1842);
assign  nx694 = ~(((nx1583) | (nx1724)) & ((src1_4) | (nx1711)));
assign  sub_result_4 = ~(((nx1569) & (~(nx1581))) | ((~(nx1569)) & (nx1581)));
assign  nx358 = ~(nx1541);
assign  nx1585 = ~((~(src2_4)) | (src1_4));
assign  nx1671 = ~(((nx350) & (src1_2)) | ((nx350) & (src2_2)) | ((src1_2) & (src2_2)));
assign  nx1674 = ~((src1_1) | (src2_1));
assign  nx1676 = ~((src1_3) | (src2_3));
assign  nx1583 = ~((src2_4) & (src1_4));
assign  nx684 = ((nx1906) & (~(nx1911))) | ((~(nx1906)) & (nx1911));
assign  nx42 = (src2_6) & ~(cycle_0) & ~(cycle_1) | (src2_4) & (cycle_0) & ~(cycle_1) | (src2_2) & ~(cycle_0) & (cycle_1) | (src2_0) & (cycle_0) & (cycle_1);
assign  nx40 = ~(nx1509);
assign  nx44 = ~((nx1537) | (nx1509));
assign  nx1868 = ~(((src1_4) & (nx114)) | ((src1_2) & (nx308)));
assign  nx1950 = ~((nx804) | ((src1_5) & (nx658)) | ((nx750) & (nx222)));
assign  nx974 = ~(((nx1611) & (nx1585)) | ((nx1611) & (src2_5)) | ((nx1585) & (src2_5)));
assign  nx1008 = ~(nx134);
assign  nx1557 = ((nx1559) & (~(nx1563))) | ((~(nx1559)) & (nx1563));
assign  des_acc_6 = ~((nx1974) & (nx1976) & (nx1978) & (nx1997));
assign  nx1000 = ~(nx204);
assign  nx1997 = ~((((nx916) | (nx900)) & (nx338)) | (nx888));
assign  nx531 = ~(((nx533) & (~(nx535))) | ((~(nx533)) & (nx535)));
assign  nx535 = ~((src1_6) & (nx42));
assign  nx536 = ~(((nx1561) | (nx1724)) & ((src1_3) | (nx1711)));
assign  nx1991 = ~((nx936) | ((src1_6) & (nx658)) | ((nx876) & (nx222)));
assign  nx1994 = ~((src1_6) | (src2_6));
assign  nx437 = ~((src1_1) & (nx72) & (mulsrc2_0));
assign  nx120 = ~(((nx484) & (~(nx487)) & (~(nx474))) | ((~(nx484)) & (nx487) & (~(nx474))) | ((~(nx484)) & (~(nx487)) & (nx474)) | ((nx484) & (nx487) & (nx474)));
assign  nx435 = ~(((nx437) & (~(nx440_mul))) | ((~(nx437)) & (nx440_mul)));
assign  divsrc2_0 = ~((nx801) | (nx826));
assign  divsrc1_1 = ~((nx861) & ((nx853) | (divsrc2_0)));
assign  nx1859 = ~(nx194);
assign  nx1862 = ((nx350) & (~(nx1541))) | ((~(nx350)) & (nx1541));
assign  nx546 = ~(nx210);
assign  divsrc1_6 = ~((nx963) & ((nx957) | (divsrc2_0)));
assign  nx1906 = ~(((nx550) & (srcCy)) | ((nx550) & (src1_3)) | ((srcCy) & (src1_3)));
assign  nx1903 = ~((nx694) | ((nx684) & (nx262)));
endmodule

module ALU ( bit_in, cycle_0, cycle_0_div, cycle_1, cycle_1_div, enable_div, enable_mul, nx10, nx102, nx110, nx114, nx12, nx128, nx136, nx1598, nx1639, nx1641, nx1696, nx1698, nx1711, nx1724, nx1763, nx1768, nx1776, nx1778, nx178, nx1782, nx18, nx1819, nx1890, nx1901, nx1922, nx1945, nx2019, nx2028, nx216, nx22, nx222, nx226, nx236, nx244, nx252, nx262, nx290, nx308, nx338, nx36, nx386, nx415, nx433, nx455, nx459, nx474, nx50, nx504, nx506, nx537, nx539, nx567, nx575, nx593, nx60, nx601, nx605, nx64, nx730, nx806, nx812, nx94, op_code_0_, op_code_1_, op_code_2_, op_code_3_, src1_0_, src1_1_, src1_2_, src1_3_, src1_4_, src1_5_, src1_6_, src1_7_, src2_0_, src2_1_, src2_2_, src2_3_, src2_4_, src2_5_, src2_6_, src2_7_, srcAc, srcCy, tmp_mul_10, tmp_mul_11, tmp_mul_12, tmp_mul_8, tmp_mul_9, tmp_rem_0, tmp_rem_1, tmp_rem_2, tmp_rem_3, tmp_rem_4, tmp_rem_5, tmp_rem_6, tmp_rem_7, desCy, des_acc_0_, des_acc_1_, des_acc_2_, des_acc_3_, des_acc_4_, des_acc_5_, des_acc_6_, des_acc_7_ );
input bit_in;
input cycle_0;
input cycle_0_div;
input cycle_1;
input cycle_1_div;
input enable_div;
input enable_mul;
input nx10;
input nx102;
input nx110;
input nx114;
input nx12;
input nx128;
input nx136;
input nx1598;
input nx1639;
input nx1641;
input nx1696;
input nx1698;
input nx1711;
input nx1724;
input nx1763;
input nx1768;
input nx1776;
input nx1778;
input nx178;
input nx1782;
input nx18;
input nx1819;
input nx1890;
input nx1901;
input nx1922;
input nx1945;
input nx2019;
input nx2028;
input nx216;
input nx22;
input nx222;
input nx226;
input nx236;
input nx244;
input nx252;
input nx262;
input nx290;
input nx308;
input nx338;
input nx36;
input nx386;
input nx415;
input nx433;
input nx455;
input nx459;
input nx474;
input nx50;
input nx504;
input nx506;
input nx537;
input nx539;
input nx567;
input nx575;
input nx593;
input nx60;
input nx601;
input nx605;
input nx64;
input nx730;
input nx806;
input nx812;
input nx94;
input op_code_0_;
input op_code_1_;
input op_code_2_;
input op_code_3_;
input src1_0_;
input src1_1_;
input src1_2_;
input src1_3_;
input src1_4_;
input src1_5_;
input src1_6_;
input src1_7_;
input src2_0_;
input src2_1_;
input src2_2_;
input src2_3_;
input src2_4_;
input src2_5_;
input src2_6_;
input src2_7_;
input srcAc;
input srcCy;
input tmp_mul_10;
input tmp_mul_11;
input tmp_mul_12;
input tmp_mul_8;
input tmp_mul_9;
input tmp_rem_0;
input tmp_rem_1;
input tmp_rem_2;
input tmp_rem_3;
input tmp_rem_4;
input tmp_rem_5;
input tmp_rem_6;
input tmp_rem_7;
output desCy;
output des_acc_0_;
output des_acc_1_;
output des_acc_2_;
output des_acc_3_;
output des_acc_4_;
output des_acc_5_;
output des_acc_6_;
output des_acc_7_;
wire des1_1_;
wire des1_2_;
wire des1_3_;
wire des1_4_;
wire des1_5_;
wire des1_6_;
wire desCy;
wire des_acc_0_;
wire des_acc_1_;
wire des_acc_2_;
wire des_acc_3_;
wire des_acc_4_;
wire des_acc_5_;
wire des_acc_6_;
wire des_acc_7_;
wire divsrc1_0;
wire divsrc1_1;
wire divsrc1_2;
wire divsrc1_3;
wire divsrc1_4;
wire divsrc1_5;
wire divsrc1_6;
wire divsrc1_7;
wire divsrc2_0;
wire divsrc2_1;
wire mulsrc1_0;
wire mulsrc1_1;
wire mulsrc1_2;
wire mulsrc1_3;
wire mulsrc1_4;
wire mulsrc1_5;
wire mulsrc1_6;
wire mulsrc1_7;
wire mulsrc2_0;
wire nx1000;
wire nx1008;
wire nx1025;
wire nx1028;
wire nx102_div;
wire nx1032;
wire nx104;
wire nx1048;
wire nx1052;
wire nx110_div;
wire nx1118;
wire nx1140;
wire nx1152;
wire nx1172;
wire nx120;
wire nx134;
wire nx146;
wire nx150;
wire nx1509;
wire nx1511;
wire nx1513;
wire nx1519;
wire nx1521;
wire nx1523;
wire nx1533;
wire nx1537;
wire nx1539;
wire nx1541;
wire nx1543;
wire nx1546;
wire nx1547;
wire nx1557;
wire nx1559;
wire nx1561;
wire nx1563;
wire nx1565;
wire nx1568;
wire nx1569;
wire nx1579;
wire nx158;
wire nx1581;
wire nx1583;
wire nx1585;
wire nx1591;
wire nx1593;
wire nx1595;
wire nx1603;
wire nx1605;
wire nx1607;
wire nx1611;
wire nx1614;
wire nx1615;
wire nx1618;
wire nx162;
wire nx1623;
wire nx1625;
wire nx1627;
wire nx1629;
wire nx1630;
wire nx1637;
wire nx1651;
wire nx1653;
wire nx1657;
wire nx1661;
wire nx1663;
wire nx1668;
wire nx1671;
wire nx1674;
wire nx1676;
wire nx1679;
wire nx168;
wire nx1681;
wire nx1685;
wire nx1687;
wire nx1689;
wire nx1706;
wire nx1714;
wire nx1718;
wire nx1730;
wire nx1733;
wire nx1736;
wire nx1739;
wire nx174;
wire nx1743;
wire nx1746;
wire nx1750;
wire nx1754;
wire nx1757;
wire nx176;
wire nx1760;
wire nx1765;
wire nx1770;
wire nx1773;
wire nx1780;
wire nx1787;
wire nx1790;
wire nx1793;
wire nx1795;
wire nx1800;
wire nx1803;
wire nx1808;
wire nx1811;
wire nx182;
wire nx1824;
wire nx1826;
wire nx1828;
wire nx1831;
wire nx1835;
wire nx1837;
wire nx1839;
wire nx1842;
wire nx1847;
wire nx1849;
wire nx1854;
wire nx1859;
wire nx1862;
wire nx1866;
wire nx1868;
wire nx1870;
wire nx1873;
wire nx1877;
wire nx188;
wire nx1880;
wire nx1882;
wire nx1887;
wire nx1894;
wire nx1896;
wire nx1898;
wire nx1903;
wire nx1906;
wire nx1911;
wire nx1914;
wire nx192;
wire nx1920;
wire nx1924;
wire nx1926;
wire nx1931;
wire nx1933;
wire nx1935;
wire nx1938;
wire nx194;
wire nx1940;
wire nx1943;
wire nx1947;
wire nx194_div;
wire nx194_mul;
wire nx1950;
wire nx1958;
wire nx1963;
wire nx1968;
wire nx1970;
wire nx1974;
wire nx1976;
wire nx1978;
wire nx1981;
wire nx1983;
wire nx1986;
wire nx1988;
wire nx1991;
wire nx1994;
wire nx1997;
wire nx200;
wire nx2000;
wire nx2002;
wire nx2004;
wire nx2006;
wire nx2013;
wire nx2016;
wire nx202;
wire nx2021;
wire nx2023;
wire nx2026;
wire nx2031;
wire nx2033;
wire nx2035;
wire nx2038;
wire nx204;
wire nx2040;
wire nx2043;
wire nx2045;
wire nx2048;
wire nx210;
wire nx214;
wire nx238;
wire nx240;
wire nx254;
wire nx258;
wire nx258_mul;
wire nx270;
wire nx298;
wire nx304;
wire nx326;
wire nx328;
wire nx330;
wire nx334;
wire nx338_mul;
wire nx342;
wire nx346;
wire nx346_div;
wire nx350;
wire nx352;
wire nx354;
wire nx358;
wire nx364;
wire nx370;
wire nx372;
wire nx374;
wire nx376;
wire nx378;
wire nx392;
wire nx396;
wire nx40;
wire nx408;
wire nx410;
wire nx410_div;
wire nx410_mul;
wire nx414;
wire nx42;
wire nx426;
wire nx428;
wire nx435;
wire nx437;
wire nx44;
wire nx440;
wire nx440_mul;
wire nx442;
wire nx442_mul;
wire nx444;
wire nx444_div;
wire nx446;
wire nx454;
wire nx458;
wire nx463;
wire nx464;
wire nx468;
wire nx471;
wire nx480;
wire nx480_div;
wire nx482;
wire nx484;
wire nx487;
wire nx489;
wire nx491;
wire nx494;
wire nx495;
wire nx498;
wire nx498_div;
wire nx500;
wire nx500_div;
wire nx502;
wire nx502_mul;
wire nx508;
wire nx510;
wire nx513;
wire nx514;
wire nx515;
wire nx516;
wire nx517;
wire nx518;
wire nx519;
wire nx520;
wire nx524;
wire nx527;
wire nx531;
wire nx533;
wire nx535;
wire nx536;
wire nx536_div;
wire nx543;
wire nx546;
wire nx550;
wire nx550_mul;
wire nx552;
wire nx552_div;
wire nx554;
wire nx554_div;
wire nx554_mul;
wire nx556;
wire nx558;
wire nx56;
wire nx561;
wire nx564;
wire nx565;
wire nx570;
wire nx572;
wire nx572_div;
wire nx579;
wire nx580;
wire nx581;
wire nx583;
wire nx588;
wire nx589;
wire nx590;
wire nx598;
wire nx603;
wire nx610;
wire nx622;
wire nx642;
wire nx648;
wire nx658;
wire nx662;
wire nx664;
wire nx680;
wire nx684;
wire nx694;
wire nx710;
wire nx714;
wire nx72;
wire nx739;
wire nx743;
wire nx744;
wire nx746;
wire nx750;
wire nx756;
wire nx76;
wire nx762;
wire nx768;
wire nx776;
wire nx78;
wire nx784;
wire nx786;
wire nx80;
wire nx801;
wire nx804;
wire nx814;
wire nx819;
wire nx821;
wire nx823;
wire nx826;
wire nx829;
wire nx832;
wire nx835;
wire nx836;
wire nx841;
wire nx843;
wire nx849;
wire nx851;
wire nx853;
wire nx855;
wire nx86;
wire nx861;
wire nx865;
wire nx868;
wire nx868_div;
wire nx870;
wire nx871;
wire nx873;
wire nx876;
wire nx879;
wire nx882;
wire nx882_div;
wire nx884;
wire nx887;
wire nx888;
wire nx890;
wire nx893;
wire nx897;
wire nx900;
wire nx901;
wire nx904;
wire nx907;
wire nx910;
wire nx910_div;
wire nx913;
wire nx915;
wire nx916;
wire nx919;
wire nx923;
wire nx926;
wire nx929;
wire nx931;
wire nx936;
wire nx937;
wire nx940;
wire nx942;
wire nx945;
wire nx946;
wire nx948;
wire nx950;
wire nx953;
wire nx957;
wire nx960;
wire nx963;
wire nx966;
wire nx974;
wire nx975;
wire nx978;
wire nx978_div;
wire nx980;
wire nx983;
wire nx986;
wire nx989;
wire nx998;
wire sub_result_0_;
wire sub_result_1_;
wire sub_result_2_;
wire sub_result_3_;
wire sub_result_4_;
wire sub_result_5_;
wire sub_result_6_;
wire sub_result_7_;
INV_X0P5B_A12TS ix1001 ( .Y(nx1000), .A(nx204) );
NAND4_X0P5A_A12TS ix1007 ( .Y(des_acc_6_), .A(nx1974), .B(nx1976), .C(nx1978), .D(nx1997) );
INV_X0P5B_A12TS ix1009 ( .Y(nx1008), .A(nx134) );
INV_X0P5B_A12TS ix1024 ( .Y(nx1025), .A(nx354) );
INV_X0P5B_A12TS ix1029 ( .Y(nx1028), .A(nx1739) );
NOR2B_X0P7M_A12TS ix1033 ( .Y(nx1032), .AN(nx910), .B(nx1739) );
OA21A1OI2_X0P5M_A12TS ix103_div ( .Y(nx102_div), .A0(src2_5_), .A1(src2_6_), .B0(nx806), .C0(src2_7_) );
AOI21_X0P5M_A12TS ix1049 ( .Y(nx1048), .A0(nx2043), .A1(nx2045), .B0(nx1778) );
AND4_X0P5M_A12TS ix105 ( .Y(nx104), .A(nx819), .B(nx821), .C(nx823), .D(nx102_div) );
OAI21_X0P5M_A12TS ix1053 ( .Y(nx1052), .A0(nx1768), .A1(nx2038), .B0(nx2040) );
XNOR2_X0P5M_A12TS ix1081 ( .Y(sub_result_7_), .A(nx1615), .B(nx1627) );
OAI222_X0P5M_A12TS ix1119 ( .Y(nx1118), .A0(src1_7_), .A1(nx1763), .B0(nx1627), .B1(nx2019), .C0(nx2021), .C1(nx2028) );
NOR2_X0P5A_A12TS ix111_div ( .Y(nx110_div), .A(src2_7_), .B(src2_6_) );
OAI222_X0P5M_A12TS ix1141 ( .Y(nx1140), .A0(nx1629), .A1(nx1763), .B0(nx2028), .B1(nx2031), .C0(nx1689), .C1(nx2019) );
XOR2_X0P5M_A12TS ix1153 ( .Y(nx1152), .A(nx1651), .B(nx1627) );
NAND4_X0P5A_A12TS ix1161 ( .Y(des_acc_7_), .A(nx2013), .B(nx2016), .C(nx2033), .D(nx2035) );
OAI21_X0P5M_A12TS ix1173 ( .Y(nx1172), .A0(nx1651), .A1(nx1689), .B0(nx1629) );
XNOR3_X0P5M_A12TS ix121 ( .Y(nx120), .A(nx484), .B(nx487), .C(nx474) );
MXIT2_X0P5M_A12TS ix135 ( .Y(nx134), .A(nx913), .B(nx989), .S0(cycle_1_div) );
CGENI_X1M_A12TS ix147 ( .CON(nx146), .A(nx484), .B(nx489), .CI(nx491) );
CGENI_X1M_A12TS ix151 ( .CON(nx150), .A(nx513), .B(nx500), .CI(nx502_mul) );
AOI21_X0P5M_A12TS ix1510 ( .Y(nx1509), .A0(src1_0_), .A1(nx1511), .B0(nx1513) );
NAND2_X0P5A_A12TS ix1512 ( .Y(nx1511), .A(src2_0_), .B(src1_0_) );
NOR2B_X0P7M_A12TS ix1514 ( .Y(nx1513), .AN(src2_0_), .B(src1_0_) );
XOR2_X0P5M_A12TS ix1520 ( .Y(nx1519), .A(nx1521), .B(nx1513) );
OAI21_X0P5M_A12TS ix1522 ( .Y(nx1521), .A0(src1_1_), .A1(src2_1_), .B0(nx1523) );
NAND2_X0P5A_A12TS ix1524 ( .Y(nx1523), .A(src2_1_), .B(src1_1_) );
INV_X0P5B_A12TS ix1534 ( .Y(nx1533), .A(src1_0_) );
INV_X0P5B_A12TS ix1538 ( .Y(nx1537), .A(srcCy) );
XNOR2_X0P5M_A12TS ix1540 ( .Y(nx1539), .A(nx1541), .B(nx454) );
OAI21_X0P5M_A12TS ix1542 ( .Y(nx1541), .A0(src1_2_), .A1(src2_2_), .B0(nx1543) );
NAND2_X0P5A_A12TS ix1544 ( .Y(nx1543), .A(src2_2_), .B(src1_2_) );
XNOR3_X0P5M_A12TS ix1547 ( .Y(nx1546), .A(nx1736), .B(srcCy), .C(nx1032) );
INV_X0P5B_A12TS ix1548 ( .Y(nx1547), .A(src1_1_) );
XOR2_X0P5M_A12TS ix1558 ( .Y(nx1557), .A(nx1559), .B(nx1563) );
OAI21_X0P5M_A12TS ix1560 ( .Y(nx1559), .A0(src1_3_), .A1(src2_3_), .B0(nx1561) );
NAND2_X0P5A_A12TS ix1562 ( .Y(nx1561), .A(src2_3_), .B(src1_3_) );
CGENI_X1M_A12TS ix1564 ( .CON(nx1563), .A(src1_2_), .B(nx454), .CI(nx1565) );
INV_X0P5B_A12TS ix1566 ( .Y(nx1565), .A(src2_2_) );
OAI31_X0P5M_A12TS ix1569 ( .Y(nx1568), .A0(nx60), .A1(bit_in), .A2(nx64), .B0(nx1750) );
XOR2_X0P5M_A12TS ix1570 ( .Y(nx1569), .A(nx580), .B(nx710) );
INV_X0P5B_A12TS ix1580 ( .Y(nx1579), .A(src1_3_) );
AOI21_X0P5M_A12TS ix1582 ( .Y(nx1581), .A0(src1_4_), .A1(nx1583), .B0(nx1585) );
NAND2_X0P5A_A12TS ix1584 ( .Y(nx1583), .A(src2_4_), .B(src1_4_) );
NOR2B_X0P7M_A12TS ix1586 ( .Y(nx1585), .AN(src2_4_), .B(src1_4_) );
MXIT2_X0P5M_A12TS ix159 ( .Y(nx158), .A(nx893), .B(nx819), .S0(cycle_1_div) );
XOR2_X0P5M_A12TS ix1592 ( .Y(nx1591), .A(nx1593), .B(nx1585) );
OAI21_X0P5M_A12TS ix1594 ( .Y(nx1593), .A0(src1_5_), .A1(src2_5_), .B0(nx1595) );
NAND2_X0P5A_A12TS ix1596 ( .Y(nx1595), .A(src2_5_), .B(src1_5_) );
XNOR2_X0P5M_A12TS ix1604 ( .Y(nx1603), .A(nx1605), .B(nx974) );
OAI21_X0P5M_A12TS ix1606 ( .Y(nx1605), .A0(src1_6_), .A1(src2_6_), .B0(nx1607) );
NAND2_X0P5A_A12TS ix1608 ( .Y(nx1607), .A(src2_6_), .B(src1_6_) );
INV_X0P5B_A12TS ix1612 ( .Y(nx1611), .A(src1_5_) );
CGENI_X1M_A12TS ix1615 ( .CON(nx1614), .A(nx1637), .B(src2_7_), .CI(nx1615) );
XNOR2_X0P5M_A12TS ix1616 ( .Y(nx1615), .A(nx978), .B(nx1623) );
NOR2_X0P5A_A12TS ix1619 ( .Y(nx1618), .A(nx1614), .B(nx1639) );
CGENI_X1M_A12TS ix1624 ( .CON(nx1623), .A(src1_6_), .B(nx974), .CI(nx1625) );
INV_X0P5B_A12TS ix1626 ( .Y(nx1625), .A(src2_6_) );
OAI21_X0P5M_A12TS ix1628 ( .Y(nx1627), .A0(src1_7_), .A1(src2_7_), .B0(nx1629) );
OAI21_X0P5M_A12TS ix163 ( .Y(nx162), .A0(nx1511), .A1(nx1763), .B0(nx1765) );
NAND2_X0P5A_A12TS ix1630 ( .Y(nx1629), .A(src2_7_), .B(src1_7_) );
OAI22_X0P5M_A12TS ix1631 ( .Y(nx1630), .A0(srcCy), .A1(nx1711), .B0(nx1714), .B1(nx1696) );
NAND4_X0P5A_A12TS ix1635 ( .Y(desCy), .A(nx1706), .B(nx1718), .C(nx1730), .D(nx1733) );
INV_X0P5B_A12TS ix1638 ( .Y(nx1637), .A(src1_7_) );
XOR2_X0P5M_A12TS ix1652 ( .Y(nx1651), .A(nx1653), .B(nx882) );
CGENI_X1M_A12TS ix1654 ( .CON(nx1653), .A(nx868), .B(src1_6_), .CI(src2_6_) );
NOR2_X0P5A_A12TS ix1658 ( .Y(nx1657), .A(src1_5_), .B(src2_5_) );
XOR2_X0P5M_A12TS ix1662 ( .Y(nx1661), .A(nx868), .B(nx1605) );
INV_X0P5B_A12TS ix1664 ( .Y(nx1663), .A(nx756) );
XNOR2_X0P5M_A12TS ix1669 ( .Y(nx1668), .A(nx622), .B(nx514) );
CGENI_X1M_A12TS ix1672 ( .CON(nx1671), .A(nx350), .B(src1_2_), .CI(src2_2_) );
NOR2_X0P5A_A12TS ix1675 ( .Y(nx1674), .A(src1_1_), .B(src2_1_) );
NOR2_X0P5A_A12TS ix1677 ( .Y(nx1676), .A(src1_3_), .B(src2_3_) );
XNOR2_X0P5M_A12TS ix1680 ( .Y(nx1679), .A(nx1671), .B(nx1559) );
INV_X0P5B_A12TS ix1682 ( .Y(nx1681), .A(nx364) );
XNOR2_X0P5M_A12TS ix1686 ( .Y(nx1685), .A(nx1511), .B(nx1521) );
INV_X0P5B_A12TS ix1688 ( .Y(nx1687), .A(nx44) );
OAI21_X0P5M_A12TS ix169 ( .Y(nx168), .A0(op_code_0_), .A1(nx1757), .B0(nx1760) );
NOR2_X0P5A_A12TS ix1690 ( .Y(nx1689), .A(src1_7_), .B(src2_7_) );
AOI211_X0P5M_A12TS ix1707 ( .Y(nx1706), .A0(src1_7_), .A1(nx102), .B0(nx1630), .C0(nx1618) );
INV_X0P5B_A12TS ix1715 ( .Y(nx1714), .A(nx1172) );
OAI31_X0P5M_A12TS ix1719 ( .Y(nx1718), .A0(nx22), .A1(nx252), .A2(nx1598), .B0(srcCy) );
AO21A1AI2_X0P5M_A12TS ix1731 ( .Y(nx1730), .A0(nx1537), .A1(nx222), .B0(nx252), .C0(bit_in) );
OA21A1OI2_X0P5M_A12TS ix1734 ( .Y(nx1733), .A0(nx1546), .A1(nx326), .B0(nx10), .C0(nx1568) );
OAI21_X0P5M_A12TS ix1737 ( .Y(nx1736), .A0(src1_6_), .A1(src1_5_), .B0(src1_7_) );
OAI31_X0P5M_A12TS ix1740 ( .Y(nx1739), .A0(src1_6_), .A1(src1_5_), .A2(src1_7_), .B0(nx1736) );
NAND2_X0P5A_A12TS ix1744 ( .Y(nx1743), .A(src1_4_), .B(nx326) );
NOR2_X0P5A_A12TS ix1747 ( .Y(nx1746), .A(src1_2_), .B(src1_1_) );
NOR2_X0P5A_A12TS ix175 ( .Y(nx174), .A(nx812), .B(nx821) );
NAND3_X0P5A_A12TS ix1751 ( .Y(nx1750), .A(nx110), .B(src1_0_), .C(nx1698) );
AOI21_X0P5M_A12TS ix1755 ( .Y(nx1754), .A0(mulsrc1_0), .A1(enable_mul), .B0(nx168) );
AOI32_X0P5M_A12TS ix1758 ( .Y(nx1757), .A0(nx1533), .A1(op_code_1_), .A2(op_code_2_), .B0(nx40), .B1(nx128) );
AO21A1AI2_X0P5M_A12TS ix1761 ( .Y(nx1760), .A0(src1_0_), .A1(nx128), .B0(nx162), .C0(op_code_0_) );
OAI21_X0P5M_A12TS ix1766 ( .Y(nx1765), .A0(nx136), .A1(nx128), .B0(src2_0_) );
INV_X0P5B_A12TS ix177 ( .Y(nx176), .A(nx950) );
AOI22_X0P5M_A12TS ix1771 ( .Y(nx1770), .A0(src1_1_), .A1(nx114), .B0(divsrc1_0), .B1(enable_div) );
AOI221_X0P5M_A12TS ix1774 ( .Y(nx1773), .A0(srcCy), .A1(nx102), .B0(sub_result_0_), .B1(nx94), .C0(nx76) );
AOI31_X0P5M_A12TS ix1781 ( .Y(nx1780), .A0(nx1641), .A1(src1_7_), .A2(nx1782), .B0(nx56) );
AOI22_X0P5M_A12TS ix1788 ( .Y(nx1787), .A0(mulsrc1_1), .A1(enable_mul), .B0(nx330), .B1(nx338) );
NOR2_X0P5A_A12TS ix1791 ( .Y(nx1790), .A(nx326), .B(srcAc) );
AOI22_X0P5M_A12TS ix1794 ( .Y(nx1793), .A0(src1_2_), .A1(nx114), .B0(divsrc1_1), .B1(enable_div) );
AOI22_X0P5M_A12TS ix1796 ( .Y(nx1795), .A0(src1_0_), .A1(nx308), .B0(sub_result_1_), .B1(nx94) );
AOI21_X0P5M_A12TS ix1801 ( .Y(nx1800), .A0(des1_1_), .A1(nx290), .B0(nx200) );
AOI222_X0P5M_A12TS ix1804 ( .Y(nx1803), .A0(nx182), .A1(nx252), .B0(src2_1_), .B1(nx244), .C0(nx258), .C1(nx262) );
XNOR2_X0P5M_A12TS ix1809 ( .Y(nx1808), .A(src1_1_), .B(srcCy) );
NAND3_X0P5A_A12TS ix181 ( .Y(des_acc_0_), .A(nx1754), .B(nx1770), .C(nx1773) );
AOI221_X0P5M_A12TS ix1812 ( .Y(nx1811), .A0(nx188), .A1(nx222), .B0(src1_1_), .B1(nx216), .C0(nx240) );
AOI22_X0P5M_A12TS ix1825 ( .Y(nx1824), .A0(mulsrc1_2), .A1(enable_mul), .B0(divsrc1_2), .B1(enable_div) );
AOI22_X0P5M_A12TS ix1827 ( .Y(nx1826), .A0(src1_3_), .A1(nx114), .B0(src1_1_), .B1(nx308) );
AOI22_X0P5M_A12TS ix1829 ( .Y(nx1828), .A0(des1_2_), .A1(nx442), .B0(sub_result_2_), .B1(nx94) );
INV_X0P5B_A12TS ix183 ( .Y(nx182), .A(nx1674) );
AOI222_X0P5M_A12TS ix1832 ( .Y(nx1831), .A0(nx352), .A1(nx252), .B0(src2_2_), .B1(nx244), .C0(nx414), .C1(nx262) );
CGENI_X1M_A12TS ix1836 ( .CON(nx1835), .A(src1_0_), .B(src1_1_), .CI(srcCy) );
XNOR2_X0P5M_A12TS ix1838 ( .Y(nx1837), .A(srcCy), .B(src1_2_) );
AOI221_X0P5M_A12TS ix1840 ( .Y(nx1839), .A0(nx358), .A1(nx222), .B0(src1_2_), .B1(nx216), .C0(nx396) );
NOR2_X0P5A_A12TS ix1843 ( .Y(nx1842), .A(src1_2_), .B(src2_2_) );
NAND4B_X0P5M_A12TS ix1848 ( .Y(nx1847), .AN(op_code_3_), .B(op_code_0_), .C(nx1790), .D(op_code_2_) );
AOI31_X0P5M_A12TS ix1850 ( .Y(nx1849), .A0(nx376), .A1(nx328), .A2(nx338), .B0(nx370) );
OAI21_X0P5M_A12TS ix1855 ( .Y(nx1854), .A0(src1_2_), .A1(src1_1_), .B0(src1_3_) );
INV_X0P5B_A12TS ix1860 ( .Y(nx1859), .A(nx194) );
XOR2_X0P5M_A12TS ix1863 ( .Y(nx1862), .A(nx350), .B(nx1541) );
AOI22_X0P5M_A12TS ix1867 ( .Y(nx1866), .A0(mulsrc1_3), .A1(enable_mul), .B0(divsrc1_3), .B1(enable_div) );
AOI22_X0P5M_A12TS ix1869 ( .Y(nx1868), .A0(src1_4_), .A1(nx114), .B0(src1_2_), .B1(nx308) );
AOI22_X0P5M_A12TS ix1871 ( .Y(nx1870), .A0(des1_3_), .A1(nx564), .B0(sub_result_3_), .B1(nx94) );
AOI222_X0P5M_A12TS ix1874 ( .Y(nx1873), .A0(nx502), .A1(nx252), .B0(src2_3_), .B1(nx244), .C0(nx554), .C1(nx262) );
CGENI_X1M_A12TS ix1878 ( .CON(nx1877), .A(nx410), .B(srcCy), .CI(src1_2_) );
XNOR2_X0P5M_A12TS ix1881 ( .Y(nx1880), .A(srcCy), .B(src1_3_) );
AOI221_X0P5M_A12TS ix1883 ( .Y(nx1882), .A0(nx508), .A1(nx222), .B0(src1_3_), .B1(nx216), .C0(nx536) );
AOI31_X0P5M_A12TS ix1888 ( .Y(nx1887), .A0(nx1854), .A1(srcAc), .A2(nx494), .B0(nx520) );
INV_X0P5B_A12TS ix189 ( .Y(nx188), .A(nx1521) );
AOI22_X0P5M_A12TS ix1895 ( .Y(nx1894), .A0(mulsrc1_4), .A1(enable_mul), .B0(divsrc1_4), .B1(enable_div) );
AOI22_X0P5M_A12TS ix1897 ( .Y(nx1896), .A0(src1_5_), .A1(nx114), .B0(src1_3_), .B1(nx308) );
AOI22_X0P5M_A12TS ix1899 ( .Y(nx1898), .A0(des1_4_), .A1(nx290), .B0(sub_result_4_), .B1(nx94) );
AOI21_X0P5M_A12TS ix1904 ( .Y(nx1903), .A0(nx684), .A1(nx262), .B0(nx694) );
CGENI_X1M_A12TS ix1907 ( .CON(nx1906), .A(nx550), .B(srcCy), .CI(src1_3_) );
XNOR2_X0P5M_A12TS ix1912 ( .Y(nx1911), .A(src1_4_), .B(srcCy) );
OA21A1OI2_X0P5M_A12TS ix1915 ( .Y(nx1914), .A0(nx664), .A1(nx252), .B0(src2_4_), .C0(nx662) );
AOI21_X0P5M_A12TS ix1921 ( .Y(nx1920), .A0(nx1537), .A1(nx244), .B0(nx216) );
INV_X0P5B_A12TS ix1925 ( .Y(nx1924), .A(src1_4_) );
AOI31_X0P5M_A12TS ix1927 ( .Y(nx1926), .A0(nx610), .A1(nx1743), .A2(nx338), .B0(nx648) );
NOR2_X0P5A_A12TS ix193 ( .Y(nx192), .A(nx812), .B(nx823) );
AOI22_X0P5M_A12TS ix1932 ( .Y(nx1931), .A0(mulsrc1_5), .A1(enable_mul), .B0(divsrc1_5), .B1(enable_div) );
AOI22_X0P5M_A12TS ix1934 ( .Y(nx1933), .A0(src1_6_), .A1(nx114), .B0(src1_4_), .B1(nx308) );
AOI22_X0P5M_A12TS ix1936 ( .Y(nx1935), .A0(des1_5_), .A1(nx290), .B0(sub_result_5_), .B1(nx94) );
XNOR2_X0P5M_A12TS ix1939 ( .Y(nx1938), .A(nx1940), .B(nx1943) );
CGENI_X1M_A12TS ix1941 ( .CON(nx1940), .A(nx680), .B(src1_4_), .CI(srcCy) );
XNOR2_X0P5M_A12TS ix1944 ( .Y(nx1943), .A(src1_5_), .B(srcCy) );
AOI22_X0P5M_A12TS ix1948 ( .Y(nx1947), .A0(nx744), .A1(nx252), .B0(src2_5_), .B1(nx664) );
NOR2_X0P5A_A12TS ix195 ( .Y(nx194), .A(nx1685), .B(nx1687) );
AOI221_X0P5M_A12TS ix1951 ( .Y(nx1950), .A0(nx750), .A1(nx222), .B0(src1_5_), .B1(nx658), .C0(nx804) );
AOI21_X0P5M_A12TS ix1959 ( .Y(nx1958), .A0(nx338), .A1(nx786), .B0(nx762) );
INV_X0P5B_A12TS ix195_div ( .Y(nx194_div), .A(nx931) );
MXIT2_X0P5M_A12TS ix195_mul ( .Y(nx194_mul), .A(nx474), .B(nx480), .S0(nx120) );
NAND2B_X0P7M_A12TS ix1964 ( .Y(nx1963), .AN(nx1743), .B(src1_5_) );
INV_X0P5B_A12TS ix1969 ( .Y(nx1968), .A(nx642) );
XNOR2_X0P5M_A12TS ix1971 ( .Y(nx1970), .A(nx1583), .B(nx1593) );
AOI22_X0P5M_A12TS ix1975 ( .Y(nx1974), .A0(mulsrc1_6), .A1(enable_mul), .B0(divsrc1_6), .B1(enable_div) );
AOI22_X0P5M_A12TS ix1977 ( .Y(nx1976), .A0(src1_7_), .A1(nx114), .B0(src1_5_), .B1(nx308) );
AOI22_X0P5M_A12TS ix1979 ( .Y(nx1978), .A0(des1_6_), .A1(nx290), .B0(sub_result_6_), .B1(nx94) );
XNOR2_X0P5M_A12TS ix1982 ( .Y(nx1981), .A(nx1983), .B(nx1986) );
CGENI_X1M_A12TS ix1984 ( .CON(nx1983), .A(nx814), .B(src1_5_), .CI(srcCy) );
XNOR2_X0P5M_A12TS ix1987 ( .Y(nx1986), .A(src1_6_), .B(srcCy) );
AOI22_X0P5M_A12TS ix1989 ( .Y(nx1988), .A0(nx870), .A1(nx252), .B0(src2_6_), .B1(nx664) );
AOI221_X0P5M_A12TS ix1992 ( .Y(nx1991), .A0(nx876), .A1(nx222), .B0(src1_6_), .B1(nx658), .C0(nx936) );
NOR2_X0P5A_A12TS ix1995 ( .Y(nx1994), .A(src1_6_), .B(src2_6_) );
OA21A1OI2_X0P5M_A12TS ix1998 ( .Y(nx1997), .A0(nx916), .A1(nx900), .B0(nx338), .C0(nx888) );
INV_X0P5B_A12TS ix2001 ( .Y(nx2000), .A(nx768) );
AOI21_X0P5M_A12TS ix2003 ( .Y(nx2002), .A0(src1_5_), .A1(src1_6_), .B0(nx2004) );
NOR2_X0P5A_A12TS ix2005 ( .Y(nx2004), .A(src1_6_), .B(src1_5_) );
INV_X0P5B_A12TS ix2007 ( .Y(nx2006), .A(nx784) );
AOI211_X0P5M_A12TS ix201 ( .Y(nx200), .A0(nx1687), .A1(nx1685), .B0(nx194), .C0(nx1696) );
NAND2_X0P5A_A12TS ix2014 ( .Y(nx2013), .A(nx1152), .B(nx50) );
MXIT2_X0P5M_A12TS ix2017 ( .Y(nx2016), .A(nx1118), .B(nx1140), .S0(op_code_0_) );
XNOR2_X0P5M_A12TS ix2022 ( .Y(nx2021), .A(nx2023), .B(nx2026) );
CGENI_X1M_A12TS ix2024 ( .CON(nx2023), .A(nx946), .B(src1_6_), .CI(srcCy) );
XNOR2_X0P5M_A12TS ix2027 ( .Y(nx2026), .A(src1_7_), .B(srcCy) );
MXIT2_X0P5M_A12TS ix203 ( .Y(nx202), .A(nx471), .B(nx506), .S0(nx510) );
MXIT2_X0P5M_A12TS ix2032 ( .Y(nx2031), .A(src1_7_), .B(src2_7_), .S0(srcCy) );
AOI22_X0P5M_A12TS ix2034 ( .Y(nx2033), .A0(mulsrc1_7), .A1(enable_mul), .B0(divsrc1_7), .B1(enable_div) );
AOI221_X0P5M_A12TS ix2036 ( .Y(nx2035), .A0(src1_7_), .A1(nx22), .B0(sub_result_7_), .B1(nx94), .C0(nx1052) );
AOI22_X0P5M_A12TS ix2039 ( .Y(nx2038), .A0(src1_0_), .A1(nx18), .B0(srcCy), .B1(nx1698) );
AOI31_X0P5M_A12TS ix2041 ( .Y(nx2040), .A0(nx1782), .A1(op_code_1_), .A2(src1_6_), .B0(nx1048) );
NAND4_X0P5A_A12TS ix2044 ( .Y(nx2043), .A(nx1854), .B(nx1537), .C(src1_7_), .D(nx2004) );
OAI211_X0P5M_A12TS ix2046 ( .Y(nx2045), .A0(nx910), .A1(nx1028), .B0(nx784), .C0(nx2048) );
INV_X0P5B_A12TS ix2049 ( .Y(nx2048), .A(nx1032) );
NOR2_X0P5A_A12TS ix205 ( .Y(nx204), .A(nx812), .B(nx913) );
CGENI_X1M_A12TS ix211 ( .CON(nx210), .A(nx527), .B(nx517), .CI(nx519) );
NOR2_X0P5A_A12TS ix215 ( .Y(nx214), .A(nx812), .B(nx893) );
NOR2B_X0P7M_A12TS ix239 ( .Y(nx238), .AN(src2_0_), .B(nx730) );
OAI22_X0P5M_A12TS ix241 ( .Y(nx240), .A0(nx1523), .A1(nx1724), .B0(src1_1_), .B1(nx1711) );
CGENI_X1M_A12TS ix255 ( .CON(nx254), .A(nx546), .B(nx533), .CI(nx535) );
AO21A1AI2_X0P5M_A12TS ix257 ( .Y(divsrc1_0), .A0(divsrc2_0), .A1(nx238), .B0(nx841), .C0(nx843) );
XNOR2_X0P5M_A12TS ix259 ( .Y(nx258), .A(src1_0_), .B(nx1808) );
CGENI_X1M_A12TS ix259_mul ( .CON(nx258_mul), .A(nx561), .B(nx552), .CI(nx554_mul) );
NAND4B_X0P5M_A12TS ix269 ( .Y(nx739), .AN(tmp_rem_0), .B(cycle_0_div), .C(cycle_1_div), .D(src2_0_) );
NAND2_X0P5A_A12TS ix271 ( .Y(des1_1_), .A(nx1803), .B(nx1811) );
XNOR2_X0P5M_A12TS ix271_div ( .Y(nx270), .A(nx739), .B(nx851) );
OAI21_X0P5M_A12TS ix275 ( .Y(divsrc1_1), .A0(nx853), .A1(divsrc2_0), .B0(nx861) );
NAND2B_X0P7M_A12TS ix299 ( .Y(nx298), .AN(nx80), .B(nx1519) );
XOR2_X0P5M_A12TS ix305 ( .Y(sub_result_1_), .A(nx80), .B(nx1519) );
MXIT2_X0P5M_A12TS ix305_mul ( .Y(nx304), .A(nx468), .B(nx539), .S0(nx543) );
XOR2_X0P5M_A12TS ix321 ( .Y(mulsrc1_1), .A(nx572), .B(nx579) );
INV_X0P5B_A12TS ix327 ( .Y(nx326), .A(nx1854) );
XNOR2_X0P5M_A12TS ix327_mul ( .Y(mulsrc1_0), .A(nx304), .B(nx556) );
INV_X0P5B_A12TS ix329 ( .Y(nx328), .A(nx1790) );
XNOR2_X0P5M_A12TS ix331 ( .Y(nx330), .A(src1_1_), .B(nx1790) );
NAND4B_X0P5M_A12TS ix335 ( .Y(nx334), .AN(tmp_rem_1), .B(src2_0_), .C(cycle_0_div), .D(cycle_1_div) );
MXIT2_X0P5M_A12TS ix339_mul ( .Y(nx338_mul), .A(nx572), .B(nx575), .S0(nx579) );
CGENI_X1M_A12TS ix343 ( .CON(nx342), .A(nx873), .B(nx897), .CI(nx214) );
NAND4_X0P5A_A12TS ix347 ( .Y(des_acc_1_), .A(nx1787), .B(nx1793), .C(nx1795), .D(nx1800) );
CGENI_X1M_A12TS ix347_div ( .CON(nx346_div), .A(nx871), .B(nx915), .CI(nx204) );
INV_X0P5B_A12TS ix347_mul ( .Y(nx346), .A(nx583) );
OAI21_X0P5M_A12TS ix351 ( .Y(nx350), .A0(nx1511), .A1(nx1674), .B0(nx1523) );
INV_X0P5B_A12TS ix353 ( .Y(nx352), .A(nx1842) );
OA21A1OI2_X0P5M_A12TS ix355 ( .Y(mulsrc1_3), .A0(nx593), .A1(nx433), .B0(nx581), .C0(nx346) );
CGENI_X1M_A12TS ix355_div ( .CON(nx354), .A(nx868_div), .B(nx953), .CI(nx176) );
INV_X0P5B_A12TS ix359 ( .Y(nx358), .A(nx1541) );
NOR2_X0P5A_A12TS ix365 ( .Y(nx364), .A(nx1862), .B(nx1859) );
NOR3_X0P5A_A12TS ix365_div ( .Y(divsrc2_1), .A(nx865), .B(nx134), .C(nx801) );
INV_X0P5B_A12TS ix367 ( .Y(mulsrc1_2), .A(nx463) );
AOI211_X0P5M_A12TS ix371 ( .Y(nx370), .A0(nx1859), .A1(nx1862), .B0(nx364), .C0(nx1696) );
AOI21_X0P5M_A12TS ix373 ( .Y(nx372), .A0(divsrc2_1), .A1(nx238), .B0(nx998) );
INV_X0P5B_A12TS ix375 ( .Y(nx374), .A(nx603) );
AO21_X0P5M_A12TS ix377 ( .Y(nx376), .A0(src1_1_), .A1(src1_2_), .B0(nx1746) );
INV_X0P5B_A12TS ix379 ( .Y(nx378), .A(nx589) );
OA21A1OI2_X0P5M_A12TS ix387 ( .Y(mulsrc1_5), .A0(nx601), .A1(nx433), .B0(nx603), .C0(nx378) );
XOR2_X0P5M_A12TS ix393 ( .Y(nx392), .A(nx835), .B(nx890) );
OA21A1OI2_X0P5M_A12TS ix395 ( .Y(mulsrc1_4), .A0(nx459), .A1(nx433), .B0(nx583), .C0(nx374) );
OAI22_X0P5M_A12TS ix397 ( .Y(nx396), .A0(nx1543), .A1(nx1724), .B0(src1_2_), .B1(nx1711) );
OAI21_X0P5M_A12TS ix397_div ( .Y(divsrc1_2), .A0(nx879), .A1(divsrc2_0), .B0(nx887) );
INV_X0P5B_A12TS ix405 ( .Y(nx746), .A(nx884) );
NOR2_X0P5A_A12TS ix409 ( .Y(nx408), .A(nx884), .B(divsrc2_1) );
INV_X0P5B_A12TS ix41 ( .Y(nx40), .A(nx1509) );
INV_X0P5B_A12TS ix411 ( .Y(nx410), .A(nx1835) );
XNOR2_X0P5M_A12TS ix411_div ( .Y(nx410_div), .A(nx334), .B(nx882_div) );
INV_X0P5B_A12TS ix411_mul ( .Y(nx410_mul), .A(nx598) );
XOR2_X0P5M_A12TS ix415 ( .Y(nx414), .A(nx1835), .B(nx1837) );
XOR2_X0P5M_A12TS ix419 ( .Y(mulsrc1_7), .A(nx598), .B(nx605) );
NAND2_X0P5A_A12TS ix423 ( .Y(des1_2_), .A(nx1831), .B(nx1839) );
OA21A1OI2_X0P5M_A12TS ix427 ( .Y(mulsrc1_6), .A0(nx455), .A1(nx433), .B0(nx589), .C0(nx410_mul) );
MXIT2_X0P5M_A12TS ix427_div ( .Y(nx426), .A(nx835), .B(nx214), .S0(nx890) );
XNOR2_X0P5M_A12TS ix429 ( .Y(nx428), .A(nx426), .B(nx910_div) );
MXT4_X0P5M_A12TS ix43 ( .Y(nx42), .A(src2_6_), .B(src2_4_), .C(src2_2_), .D(src2_0_), .S0(cycle_0), .S1(cycle_1) );
OAI21_X0P5M_A12TS ix433_div ( .Y(divsrc1_3), .A0(nx901), .A1(divsrc2_0), .B0(nx907) );
XNOR2_X0P5M_A12TS ix436 ( .Y(nx435), .A(nx437), .B(nx440_mul) );
NAND3_X0P5A_A12TS ix438 ( .Y(nx437), .A(src1_1_), .B(nx72), .C(mulsrc2_0) );
OAI21_X0P5M_A12TS ix441 ( .Y(nx440), .A0(op_code_0_), .A1(nx12), .B0(nx1847) );
XNOR2_X0P5M_A12TS ix441_mul ( .Y(nx440_mul), .A(nx442_mul), .B(nx444) );
NAND2B_X0P7M_A12TS ix443 ( .Y(nx442), .AN(nx440), .B(nx1819) );
NAND2_X0P5A_A12TS ix443_mul ( .Y(nx442_mul), .A(src1_1_), .B(nx72) );
NAND2_X0P5A_A12TS ix445 ( .Y(nx444), .A(src1_2_), .B(nx42) );
NOR2_X0P5A_A12TS ix445_div ( .Y(nx444_div), .A(nx897), .B(divsrc2_1) );
XOR2_X0P5M_A12TS ix447 ( .Y(nx446), .A(nx873), .B(nx904) );
NOR2_X0P5A_A12TS ix45 ( .Y(nx44), .A(nx1537), .B(nx1509) );
CGENI_X1M_A12TS ix455 ( .CON(nx454), .A(nx1547), .B(nx1513), .CI(src2_1_) );
NAND2B_X0P7M_A12TS ix459 ( .Y(nx458), .AN(nx298), .B(nx1539) );
AND2_X0P5M_A12TS ix45_mul ( .Y(mulsrc2_0), .A(src1_0_), .B(nx42) );
AO21A1AI2_X0P5M_A12TS ix464 ( .Y(nx463), .A0(tmp_mul_8), .A1(nx386), .B0(nx338_mul), .C0(nx581) );
XOR2_X0P5M_A12TS ix465 ( .Y(sub_result_2_), .A(nx298), .B(nx1539) );
XOR2_X0P5M_A12TS ix465_div ( .Y(nx464), .A(nx832), .B(nx929) );
MXIT2_X0P5M_A12TS ix469 ( .Y(nx468), .A(nx202), .B(nx226), .S0(nx524) );
OAI21_X0P5M_A12TS ix469_div ( .Y(divsrc1_4), .A0(nx919), .A1(divsrc2_0), .B0(nx926) );
MXIT2_X0P5M_A12TS ix472 ( .Y(nx471), .A(nx194_mul), .B(nx178), .S0(nx495) );
INV_X0P5B_A12TS ix481 ( .Y(nx480), .A(nx86) );
NOR2_X0P5A_A12TS ix481_div ( .Y(nx480_div), .A(nx915), .B(divsrc2_1) );
XNOR2_X0P5M_A12TS ix483 ( .Y(nx482), .A(nx342), .B(nx923) );
OAI211_X0P5M_A12TS ix485 ( .Y(nx484), .A0(mulsrc2_0), .A1(nx78), .B0(src1_1_), .C0(nx72) );
NAND4_X0P5A_A12TS ix487 ( .Y(des_acc_2_), .A(nx1824), .B(nx1826), .C(nx1828), .D(nx1849) );
XNOR2_X0P5M_A12TS ix488 ( .Y(nx487), .A(nx489), .B(nx491) );
NAND2_X0P5A_A12TS ix490 ( .Y(nx489), .A(src1_2_), .B(nx72) );
NAND2_X0P5A_A12TS ix492 ( .Y(nx491), .A(src1_3_), .B(nx42) );
AOI21_X0P5M_A12TS ix495 ( .Y(nx494), .A0(nx1746), .A1(nx1579), .B0(nx1890) );
XNOR3_X0P5M_A12TS ix496 ( .Y(nx495), .A(nx146), .B(nx498), .C(nx504) );
XNOR2_X0P5M_A12TS ix499 ( .Y(nx498), .A(nx500), .B(nx502_mul) );
MXIT2_X0P5M_A12TS ix499_div ( .Y(nx498_div), .A(nx832), .B(nx194_div), .S0(nx929) );
NAND2_X0P5A_A12TS ix501 ( .Y(nx500), .A(src1_3_), .B(nx72) );
XNOR2_X0P5M_A12TS ix501_div ( .Y(nx500_div), .A(nx498_div), .B(nx948) );
INV_X0P5B_A12TS ix503 ( .Y(nx502), .A(nx1676) );
NAND2_X0P5A_A12TS ix503_mul ( .Y(nx502_mul), .A(src1_4_), .B(nx42) );
OAI21_X0P5M_A12TS ix505_div ( .Y(divsrc1_5), .A0(nx937), .A1(divsrc2_0), .B0(nx945) );
INV_X0P5B_A12TS ix509 ( .Y(nx508), .A(nx1559) );
XNOR3_X0P5M_A12TS ix511 ( .Y(nx510), .A(nx150), .B(nx515), .C(nx506) );
INV_X0P5B_A12TS ix513 ( .Y(nx743), .A(nx942) );
INV_X0P5B_A12TS ix514 ( .Y(nx513), .A(nx146) );
NOR2_X0P5A_A12TS ix515 ( .Y(nx514), .A(nx1679), .B(nx1681) );
XNOR2_X0P5M_A12TS ix516 ( .Y(nx515), .A(nx517), .B(nx519) );
NOR2_X0P5A_A12TS ix517 ( .Y(nx516), .A(nx942), .B(divsrc2_1) );
NAND2_X0P5A_A12TS ix518 ( .Y(nx517), .A(src1_4_), .B(nx72) );
XNOR2_X0P5M_A12TS ix519 ( .Y(nx518), .A(nx346_div), .B(nx940) );
NAND2_X0P5A_A12TS ix520 ( .Y(nx519), .A(src1_5_), .B(nx42) );
AOI211_X0P5M_A12TS ix521 ( .Y(nx520), .A0(nx1681), .A1(nx1679), .B0(nx514), .C0(nx1696) );
XNOR3_X0P5M_A12TS ix525 ( .Y(nx524), .A(nx210), .B(nx531), .C(nx537) );
INV_X0P5B_A12TS ix528 ( .Y(nx527), .A(nx150) );
XNOR2_X0P5M_A12TS ix532 ( .Y(nx531), .A(nx533), .B(nx535) );
NAND2_X0P5A_A12TS ix534 ( .Y(nx533), .A(src1_5_), .B(nx72) );
NAND2_X0P5A_A12TS ix536 ( .Y(nx535), .A(src1_6_), .B(nx42) );
OAI22_X0P5M_A12TS ix537 ( .Y(nx536), .A0(nx1561), .A1(nx1724), .B0(src1_3_), .B1(nx1711) );
XOR2_X0P5M_A12TS ix537_div ( .Y(nx536_div), .A(nx829), .B(nx966) );
OAI21_X0P5M_A12TS ix541 ( .Y(divsrc1_6), .A0(nx957), .A1(divsrc2_0), .B0(nx963) );
XNOR3_X0P5M_A12TS ix544 ( .Y(nx543), .A(nx254), .B(nx550_mul), .C(nx539) );
INV_X0P5B_A12TS ix547 ( .Y(nx546), .A(nx210) );
INV_X0P5B_A12TS ix551 ( .Y(nx550), .A(nx1877) );
XNOR2_X0P5M_A12TS ix551_mul ( .Y(nx550_mul), .A(nx552), .B(nx554_mul) );
NAND2_X0P5A_A12TS ix553 ( .Y(nx552), .A(src1_6_), .B(nx72) );
NOR2_X0P5A_A12TS ix553_div ( .Y(nx552_div), .A(nx953), .B(divsrc2_1) );
XOR2_X0P5M_A12TS ix555 ( .Y(nx554), .A(nx1877), .B(nx1880) );
XOR2_X0P5M_A12TS ix555_div ( .Y(nx554_div), .A(nx868_div), .B(nx960) );
NAND2_X0P5A_A12TS ix555_mul ( .Y(nx554_mul), .A(src1_7_), .B(nx42) );
XNOR2_X0P5M_A12TS ix557 ( .Y(nx556), .A(nx558), .B(nx567) );
AO21A1AI2_X0P5M_A12TS ix559 ( .Y(nx558), .A0(src1_7_), .A1(nx72), .B0(nx258_mul), .C0(nx565) );
INV_X0P5B_A12TS ix562 ( .Y(nx561), .A(nx254) );
NAND2_X0P5A_A12TS ix563 ( .Y(des1_3_), .A(nx1873), .B(nx1882) );
NAND2B_X0P7M_A12TS ix565 ( .Y(nx564), .AN(nx440), .B(nx1819) );
NAND3_X0P5A_A12TS ix566 ( .Y(nx565), .A(nx258_mul), .B(src1_7_), .C(nx72) );
AOI211_X0P5M_A12TS ix57 ( .Y(nx56), .A0(nx1509), .A1(nx1537), .B0(nx44), .C0(nx1696) );
MXIT2_X0P5M_A12TS ix571 ( .Y(nx570), .A(nx829), .B(nx158), .S0(nx966) );
MXIT2_X0P5M_A12TS ix573 ( .Y(nx572), .A(nx304), .B(nx236), .S0(nx556) );
XNOR2_X0P5M_A12TS ix573_div ( .Y(nx572_div), .A(nx570), .B(nx986) );
OAI21_X0P5M_A12TS ix577 ( .Y(divsrc1_7), .A0(nx975), .A1(divsrc2_0), .B0(nx983) );
XNOR2_X0P5M_A12TS ix580 ( .Y(nx579), .A(nx565), .B(nx575) );
NAND2B_X0P7M_A12TS ix581 ( .Y(nx580), .AN(nx458), .B(nx1557) );
NAND3_X0P5A_A12TS ix582 ( .Y(nx581), .A(nx386), .B(tmp_mul_8), .C(nx338_mul) );
NAND3B_X0P5M_A12TS ix584 ( .Y(nx583), .AN(nx581), .B(nx386), .C(tmp_mul_9) );
XOR2_X0P5M_A12TS ix587 ( .Y(sub_result_3_), .A(nx458), .B(nx1557) );
NOR2_X0P5A_A12TS ix589 ( .Y(nx588), .A(nx980), .B(divsrc2_1) );
NAND3_X0P5A_A12TS ix590 ( .Y(nx589), .A(nx386), .B(tmp_mul_11), .C(nx374) );
XNOR2_X0P5M_A12TS ix591 ( .Y(nx590), .A(nx354), .B(nx978_div) );
NAND3_X0P5A_A12TS ix599 ( .Y(nx598), .A(nx386), .B(tmp_mul_12), .C(nx378) );
NAND3_X0P5A_A12TS ix604 ( .Y(nx603), .A(nx386), .B(tmp_mul_10), .C(nx346) );
NAND4_X0P5A_A12TS ix609 ( .Y(des_acc_3_), .A(nx1866), .B(nx1868), .C(nx1870), .D(nx1887) );
NOR2_X0P5A_A12TS ix609_div ( .Y(divsrc2_0), .A(nx801), .B(nx826) );
NAND2B_X0P7M_A12TS ix611 ( .Y(nx610), .AN(src1_4_), .B(nx1854) );
OAI21_X0P5M_A12TS ix623 ( .Y(nx622), .A0(nx1671), .A1(nx1676), .B0(nx1561) );
NOR2_X0P5A_A12TS ix643 ( .Y(nx642), .A(nx1668), .B(nx1581) );
AOI211_X0P5M_A12TS ix649 ( .Y(nx648), .A0(nx1581), .A1(nx1668), .B0(nx642), .C0(nx1696) );
INV_X0P5B_A12TS ix659 ( .Y(nx658), .A(nx1920) );
AOI21_X0P5M_A12TS ix663 ( .Y(nx662), .A0(nx1920), .A1(nx1922), .B0(nx1924) );
AND2_X0P5M_A12TS ix665 ( .Y(nx664), .A(srcCy), .B(nx244) );
INV_X0P5B_A12TS ix681 ( .Y(nx680), .A(nx1906) );
XOR2_X0P5M_A12TS ix685 ( .Y(nx684), .A(nx1906), .B(nx1911) );
OAI22_X0P5M_A12TS ix695 ( .Y(nx694), .A0(nx1583), .A1(nx1724), .B0(src1_4_), .B1(nx1711) );
OAI211_X1M_A12TS ix699 ( .Y(des1_4_), .A0(nx1581), .A1(nx1901), .B0(nx1903), .C0(nx1914) );
CGENI_X1M_A12TS ix711 ( .CON(nx710), .A(nx1579), .B(nx1563), .CI(src2_3_) );
NAND2_X0P5A_A12TS ix715 ( .Y(nx714), .A(nx1581), .B(nx1569) );
XNOR2_X0P5M_A12TS ix721 ( .Y(sub_result_4_), .A(nx1569), .B(nx1581) );
MXT4_X0P5M_A12TS ix73 ( .Y(nx72), .A(src2_7_), .B(src2_5_), .C(src2_3_), .D(src2_1_), .S0(cycle_0), .S1(cycle_1) );
NAND4_X0P5A_A12TS ix743 ( .Y(des_acc_4_), .A(nx1894), .B(nx1896), .C(nx1898), .D(nx1926) );
INV_X0P5B_A12TS ix745 ( .Y(nx744), .A(nx1657) );
INV_X0P5B_A12TS ix751 ( .Y(nx750), .A(nx1593) );
NOR2_X0P5A_A12TS ix757 ( .Y(nx756), .A(nx1970), .B(nx1968) );
AOI211_X0P5M_A12TS ix763 ( .Y(nx762), .A0(nx1968), .A1(nx1970), .B0(nx756), .C0(nx1696) );
NOR2_X0P5A_A12TS ix769 ( .Y(nx768), .A(src1_5_), .B(nx1743) );
AO21A1AI2_X0P5M_A12TS ix77 ( .Y(nx76), .A0(nx1776), .A1(nx1778), .B0(nx1533), .C0(nx1780) );
OAI21_X0P5M_A12TS ix777 ( .Y(nx776), .A0(src1_5_), .A1(nx768), .B0(nx1963) );
NAND3_X0P5A_A12TS ix785 ( .Y(nx784), .A(nx1854), .B(nx1537), .C(nx1736) );
XNOR2_X0P5M_A12TS ix787 ( .Y(nx786), .A(nx776), .B(nx784) );
INV_X0P5B_A12TS ix79 ( .Y(nx78), .A(nx444) );
OA21A1OI2_X0P5M_A12TS ix802 ( .Y(nx801), .A0(nx110_div), .A1(cycle_0_div), .B0(cycle_1_div), .C0(nx104) );
OAI22_X0P5M_A12TS ix805 ( .Y(nx804), .A0(nx1595), .A1(nx1724), .B0(src1_5_), .B1(nx1711) );
NAND2_X0P5A_A12TS ix81 ( .Y(nx80), .A(nx1509), .B(srcCy) );
INV_X0P5B_A12TS ix815 ( .Y(nx814), .A(nx1940) );
MXIT2_X0P5M_A12TS ix820 ( .Y(nx819), .A(src2_4_), .B(src2_6_), .S0(cycle_0_div) );
MXIT2_X0P5M_A12TS ix822 ( .Y(nx821), .A(src2_3_), .B(src2_5_), .S0(cycle_0_div) );
MXIT2_X0P5M_A12TS ix824 ( .Y(nx823), .A(src2_2_), .B(src2_4_), .S0(cycle_0_div) );
MXIT2_X0P5M_A12TS ix827 ( .Y(nx826), .A(nx570), .B(nx1008), .S0(nx986) );
MXIT2_X0P5M_A12TS ix830 ( .Y(nx829), .A(nx498_div), .B(nx950), .S0(nx948) );
OAI211_X1M_A12TS ix831 ( .Y(des1_5_), .A0(nx1938), .A1(nx1945), .B0(nx1947), .C0(nx1950) );
MXIT2_X0P5M_A12TS ix833 ( .Y(nx832), .A(nx426), .B(nx1000), .S0(nx910_div) );
MXIT2_X0P5M_A12TS ix836 ( .Y(nx835), .A(nx739), .B(nx849), .S0(nx851) );
NAND2B_X0P7M_A12TS ix837 ( .Y(nx836), .AN(nx714), .B(nx1591) );
AOI32_X0P5M_A12TS ix842 ( .Y(nx841), .A0(src1_0_), .A1(nx806), .A2(nx812), .B0(tmp_rem_0), .B1(nx36) );
XOR2_X0P5M_A12TS ix843 ( .Y(sub_result_5_), .A(nx714), .B(nx1591) );
NAND2B_X0P7M_A12TS ix844 ( .Y(nx843), .AN(nx739), .B(divsrc2_0) );
NAND3_X0P5A_A12TS ix850 ( .Y(nx849), .A(src2_1_), .B(cycle_0_div), .C(cycle_1_div) );
XOR2_X0P5M_A12TS ix852 ( .Y(nx851), .A(nx849), .B(nx853) );
AOI21_X0P5M_A12TS ix854 ( .Y(nx853), .A0(nx855), .A1(divsrc2_1), .B0(nx372) );
INV_X0P5B_A12TS ix856 ( .Y(nx855), .A(nx334) );
NAND2_X0P5A_A12TS ix862 ( .Y(nx861), .A(divsrc2_0), .B(nx270) );
NAND4_X0P5A_A12TS ix865 ( .Y(des_acc_5_), .A(nx1931), .B(nx1933), .C(nx1935), .D(nx1958) );
CGEN_X1M_A12TS ix866 ( .CO(nx865), .A(nx1025), .B(nx980), .CI(nx158) );
OAI21_X0P5M_A12TS ix869 ( .Y(nx868), .A0(nx1583), .A1(nx1657), .B0(nx1595) );
CGENI_X1M_A12TS ix869_div ( .CON(nx868_div), .A(nx346_div), .B(nx743), .CI(nx931) );
NOR3_X0P5A_A12TS ix87 ( .Y(nx86), .A(nx433), .B(nx415), .C(nx435) );
INV_X0P5B_A12TS ix871 ( .Y(nx870), .A(nx1994) );
INV_X0P5B_A12TS ix872 ( .Y(nx871), .A(nx342) );
CGENI_X1M_A12TS ix874 ( .CON(nx873), .A(nx334), .B(nx746), .CI(nx849) );
INV_X0P5B_A12TS ix877 ( .Y(nx876), .A(nx1605) );
AOI21_X0P5M_A12TS ix880 ( .Y(nx879), .A0(divsrc2_1), .A1(nx410_div), .B0(nx408) );
NOR2_X0P5A_A12TS ix883 ( .Y(nx882), .A(nx1661), .B(nx1663) );
XOR2_X0P5M_A12TS ix883_div ( .Y(nx882_div), .A(nx884), .B(nx849) );
AOI32_X0P5M_A12TS ix885 ( .Y(nx884), .A0(src1_2_), .A1(nx806), .A2(nx812), .B0(tmp_rem_2), .B1(nx36) );
NAND2_X0P5A_A12TS ix888 ( .Y(nx887), .A(divsrc2_0), .B(nx392) );
AOI211_X0P5M_A12TS ix889 ( .Y(nx888), .A0(nx1663), .A1(nx1661), .B0(nx882), .C0(nx1696) );
OAI21_X0P5M_A12TS ix89 ( .Y(sub_result_0_), .A0(srcCy), .A1(nx1509), .B0(nx80) );
XNOR2_X0P5M_A12TS ix891 ( .Y(nx890), .A(nx214), .B(nx879) );
MXIT2_X0P5M_A12TS ix894 ( .Y(nx893), .A(src2_0_), .B(src2_2_), .S0(cycle_0_div) );
AOI32_X0P5M_A12TS ix898 ( .Y(nx897), .A0(src1_3_), .A1(nx806), .A2(nx812), .B0(tmp_rem_3), .B1(nx36) );
AND4_X0P5M_A12TS ix901 ( .Y(nx900), .A(nx1854), .B(src1_6_), .C(nx1537), .D(nx1736) );
AOI21_X0P5M_A12TS ix902 ( .Y(nx901), .A0(divsrc2_1), .A1(nx446), .B0(nx444_div) );
XNOR2_X0P5M_A12TS ix905 ( .Y(nx904), .A(nx897), .B(nx214) );
NAND2_X0P5A_A12TS ix908 ( .Y(nx907), .A(divsrc2_0), .B(nx428) );
NOR3_X0P5A_A12TS ix911 ( .Y(nx910), .A(src1_5_), .B(src1_6_), .C(nx1743) );
XNOR2_X0P5M_A12TS ix911_div ( .Y(nx910_div), .A(nx204), .B(nx901) );
MXIT2_X0P5M_A12TS ix914 ( .Y(nx913), .A(src2_1_), .B(src2_3_), .S0(cycle_0_div) );
AOI32_X0P5M_A12TS ix916 ( .Y(nx915), .A0(src1_4_), .A1(nx806), .A2(nx812), .B0(tmp_rem_4), .B1(nx36) );
AOI211_X0P5M_A12TS ix917 ( .Y(nx916), .A0(nx2000), .A1(nx2002), .B0(nx2006), .C0(nx910) );
AOI21_X0P5M_A12TS ix920 ( .Y(nx919), .A0(divsrc2_1), .A1(nx482), .B0(nx480_div) );
XNOR2_X0P5M_A12TS ix924 ( .Y(nx923), .A(nx915), .B(nx204) );
NAND2_X0P5A_A12TS ix927 ( .Y(nx926), .A(divsrc2_0), .B(nx464) );
XOR2_X0P5M_A12TS ix930 ( .Y(nx929), .A(nx931), .B(nx919) );
AOI31_X0P5M_A12TS ix932 ( .Y(nx931), .A0(cycle_0_div), .A1(src2_0_), .A2(nx812), .B0(nx192) );
OAI22_X0P5M_A12TS ix937 ( .Y(nx936), .A0(nx1607), .A1(nx1724), .B0(src1_6_), .B1(nx1711) );
AOI21_X0P5M_A12TS ix938 ( .Y(nx937), .A0(divsrc2_1), .A1(nx518), .B0(nx516) );
XOR2_X0P5M_A12TS ix941 ( .Y(nx940), .A(nx942), .B(nx931) );
AOI32_X0P5M_A12TS ix943 ( .Y(nx942), .A0(src1_5_), .A1(nx806), .A2(nx812), .B0(tmp_rem_5), .B1(nx36) );
NAND2_X0P5A_A12TS ix946 ( .Y(nx945), .A(divsrc2_0), .B(nx500_div) );
INV_X0P5B_A12TS ix947 ( .Y(nx946), .A(nx1983) );
XOR2_X0P5M_A12TS ix949 ( .Y(nx948), .A(nx950), .B(nx937) );
AOI31_X0P5M_A12TS ix951 ( .Y(nx950), .A0(cycle_0_div), .A1(src2_1_), .A2(nx812), .B0(nx174) );
AOI32_X0P5M_A12TS ix954 ( .Y(nx953), .A0(src1_6_), .A1(nx806), .A2(nx812), .B0(tmp_rem_6), .B1(nx36) );
AOI21_X0P5M_A12TS ix958 ( .Y(nx957), .A0(divsrc2_1), .A1(nx554_div), .B0(nx552_div) );
XOR2_X0P5M_A12TS ix961 ( .Y(nx960), .A(nx953), .B(nx950) );
OAI211_X1M_A12TS ix963 ( .Y(des1_6_), .A0(nx1981), .A1(nx1945), .B0(nx1988), .C0(nx1991) );
NAND2_X0P5A_A12TS ix964 ( .Y(nx963), .A(divsrc2_0), .B(nx536_div) );
XNOR2_X0P5M_A12TS ix967 ( .Y(nx966), .A(nx158), .B(nx957) );
CGENI_X1M_A12TS ix975 ( .CON(nx974), .A(nx1611), .B(nx1585), .CI(src2_5_) );
AOI21_X0P5M_A12TS ix976 ( .Y(nx975), .A0(nx590), .A1(divsrc2_1), .B0(nx588) );
NAND2B_X0P7M_A12TS ix979 ( .Y(nx978), .AN(nx836), .B(nx1603) );
XNOR2_X0P5M_A12TS ix979_div ( .Y(nx978_div), .A(nx980), .B(nx158) );
AOI32_X0P5M_A12TS ix981 ( .Y(nx980), .A0(src1_7_), .A1(nx806), .A2(nx812), .B0(tmp_rem_7), .B1(nx36) );
NAND2_X0P5A_A12TS ix984 ( .Y(nx983), .A(nx572_div), .B(divsrc2_0) );
XOR2_X0P5M_A12TS ix985 ( .Y(sub_result_6_), .A(nx836), .B(nx1603) );
XNOR2_X0P5M_A12TS ix987 ( .Y(nx986), .A(nx134), .B(nx975) );
MXIT2_X0P5M_A12TS ix990 ( .Y(nx989), .A(src2_5_), .B(src2_7_), .S0(cycle_0_div) );
AOI32_X0P5M_A12TS ix999 ( .Y(nx998), .A0(src1_1_), .A1(nx806), .A2(nx812), .B0(tmp_rem_1), .B1(nx36) );
endmodule

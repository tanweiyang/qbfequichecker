module ALU ( nx474, des_acc_7_ );

input nx474;
output des_acc_7_;
wire nx471; 

assign  des_acc_7_ = nx471 & nx474;

endmodule
